module test(a15, a14, a13, a12, a11, a10, a9, a8, a7, a6, a5, a4, a3,
     a2, a1, a0, b15, b14, b13, b12, b11, b10, b9, b8, b7, b6, b5, b4,
     b3, b2, b1, b0, o15, o14, o13, o12, o11, o10, o9, o8, o7, o6, o5,
     o4, o3, o2, o1, o0);
  input a15, a14, a13, a12, a11, a10, a9, a8, a7, a6, a5, a4, a3, a2,
       a1, a0, b15, b14, b13, b12, b11, b10, b9, b8, b7, b6, b5, b4,
       b3, b2, b1, b0;
  output o15, o14, o13, o12, o11, o10, o9, o8, o7, o6, o5, o4, o3, o2,
       o1, o0;
  wire a15, a14, a13, a12, a11, a10, a9, a8, a7, a6, a5, a4, a3, a2,
       a1, a0, b15, b14, b13, b12, b11, b10, b9, b8, b7, b6, b5, b4,
       b3, b2, b1, b0;
  wire o15, o14, o13, o12, o11, o10, o9, o8, o7, o6, o5, o4, o3, o2,
       o1, o0;
  wire n_9315, n_9316, n_9317, n_9318, n_9319, n_9320, n_9321, n_9322;
  wire n_9323, n_9324, n_9325, n_9326, n_9327, n_9328, n_9329, n_9330;
  wire n_9331, n_9332, n_9333, n_9334, n_9335, n_9337, n_9338, n_9339;
  wire n_9340, n_9341, n_9342, n_9343, n_9344, n_9345, n_9346, n_9347;
  wire n_9348, n_9349, n_9350, n_9351, n_9352, n_9353, n_9354, n_9355;
  wire n_9356, n_9357, n_9358, n_9359, n_9360, n_9361, n_9362, n_9363;
  wire n_9364, n_9365, n_9366, n_9367, n_9368, n_9369, n_9370, n_9371;
  wire n_9372, n_9373, n_9374, n_9375, n_9376, n_9377, n_9378, n_9379;
  wire n_9380, n_9381, n_9382, n_9383, n_9384, n_9385, n_9386, n_9387;
  wire n_9389, n_9390, n_9391, n_9392, n_9393, n_9394, n_9396, n_9397;
  wire n_9398, n_9399, n_9400, n_9401, n_9402, n_9403, n_9404, n_9405;
  wire n_9406, n_9407, n_9408, n_9409, n_9410, n_9411, n_9413, n_9414;
  wire n_9415, n_9416, n_9417, n_9418, n_9419, n_9420, n_9421, n_9422;
  wire n_9423, n_9424, n_9425, n_9426, n_9428, n_9429, n_9430, n_9431;
  wire n_9432, n_9433, n_9434, n_9435, n_9436, n_9437, n_9438, n_9439;
  wire n_9440, n_9441, n_9442, n_9443, n_9444, n_9445, n_9446, n_9447;
  wire n_9448, n_9449, n_9451, n_9452, n_9453, n_9454, n_9455, n_9456;
  wire n_9457, n_9458, n_9459, n_9460, n_9461, n_9462, n_9463, n_9464;
  wire n_9465, n_9466, n_9467, n_9468, n_9469, n_9470, n_9471, n_9472;
  wire n_9473, n_9474, n_9475, n_9476, n_9477, n_9478, n_9479, n_9480;
  wire n_9481, n_9482, n_9483, n_9484, n_9485, n_9486, n_9487, n_9488;
  wire n_9489, n_9490, n_9491, n_9492, n_9493, n_9494, n_9495, n_9496;
  wire n_9497, n_9498, n_9499, n_9500, n_9501, n_9503, n_9504, n_9505;
  wire n_9506, n_9507, n_9508, n_9509, n_9510, n_9511, n_9512, n_9513;
  wire n_9514, n_9515, n_9516, n_9517, n_9518, n_9519, n_9520, n_9521;
  wire n_9522, n_9523, n_9524, n_9525, n_9526, n_9527, n_9528, n_9529;
  wire n_9530, n_9531, n_9532, n_9533, n_9534, n_9535, n_9536, n_9537;
  wire n_9538, n_9540, n_9541, n_9542, n_9543, n_9544, n_9545, n_9546;
  wire n_9547, n_9548, n_9549, n_9550, n_9551, n_9552, n_9553, n_9554;
  wire n_9555, n_9556, n_9557, n_9558, n_9559, n_9560, n_9561, n_9562;
  wire n_9563, n_9564, n_9565, n_9566, n_9567, n_9568, n_9570, n_9572;
  wire n_9573, n_9574, n_9575, n_9576, n_9577, n_9578, n_9579, n_9580;
  wire n_9581, n_9582, n_9583, n_9584, n_9585, n_9586, n_9587, n_9588;
  wire n_9589, n_9590, n_9591, n_9592, n_9593, n_9594, n_9595, n_9596;
  wire n_9597, n_9598, n_9599, n_9600, n_9601, n_9602, n_9603, n_9604;
  wire n_9605, n_9606, n_9607, n_9608, n_9609, n_9610, n_9611, n_9612;
  wire n_9613, n_9614, n_9615, n_9616, n_9617, n_9618, n_9619, n_9620;
  wire n_9621, n_9622, n_9623, n_9624, n_9625, n_9626, n_9627, n_9628;
  wire n_9629, n_9630, n_9631, n_9632, n_9633, n_9634, n_9635, n_9636;
  wire n_9637, n_9638, n_9639, n_9640, n_9641, n_9642, n_9643, n_9644;
  wire n_9645, n_9646, n_9647, n_9648, n_9649, n_9650, n_9652, n_9653;
  wire n_9654, n_9655, n_9656, n_9657, n_9658, n_9659, n_9660, n_9661;
  wire n_9662, n_9663, n_9664, n_9665, n_9666, n_9667, n_9668, n_9669;
  wire n_9670, n_9671, n_9672, n_9673, n_9674, n_9675, n_9676, n_9677;
  wire n_9678, n_9679, n_9680, n_9681, n_9682, n_9683, n_9684, n_9685;
  wire n_9686, n_9687, n_9688, n_9689, n_9690, n_9691, n_9692, n_9693;
  wire n_9694, n_9695, n_9696, n_9697, n_9698, n_9699, n_9700, n_9701;
  wire n_9702, n_9703, n_9704, n_9705, n_9706, n_9707, n_9708, n_9709;
  wire n_9710, n_9711, n_9712, n_9713, n_9714, n_9715, n_9716, n_9717;
  wire n_9718, n_9719, n_9720, n_9721, n_9722, n_9723, n_9724, n_9725;
  wire n_9726, n_9727, n_9728, n_9729, n_9730, n_9731, n_9732, n_9733;
  wire n_9734, n_9735, n_9736, n_9737, n_9738, n_9739, n_9740, n_9741;
  wire n_9742, n_9743, n_9744, n_9745, n_9746, n_9747, n_9748, n_9749;
  wire n_9750, n_9751, n_9760, n_9761, n_9762, n_9763, n_9764, n_9765;
  wire n_9766, n_9767, n_9768, n_9769, n_9770, n_9771, n_9772, n_9773;
  wire n_9774, n_9775, n_9776, n_9777, n_9778, n_9779, n_9780, n_9781;
  wire n_9782, n_9783, n_9784, n_9785, n_9786, n_9787, n_9788, n_9792;
  wire n_9799, n_9800, n_9801, n_9802, n_9807, n_9808, n_9809, n_9812;
  wire n_9815, n_9816, n_9817, n_9818, n_9822, n_9826, n_9827, n_9828;
  wire n_9831, n_9838, n_9839, n_9841, n_9843, n_9846, n_9848, n_9850;
  wire n_9851, n_9852, n_9853, n_9856, n_9861, n_9862, n_9863, n_9864;
  wire n_9866, n_9867, n_9868, n_9869, n_9871, n_9873, n_9874, n_9875;
  wire n_9879, n_9880, n_9881, n_9884, n_9886, n_9887, n_9889, n_9894;
  wire n_9895, n_9896, n_9897, n_9898, n_9899, n_9900, n_9901, n_9902;
  wire n_9903, n_9904, n_9905, n_9906, n_9907, n_9908, n_9909, n_9910;
  wire n_9912, n_9914, n_9915, n_9916, n_9917, n_9918, n_9919, n_9920;
  wire n_9921, n_9922, n_9924, n_9925, n_9927, n_9928, n_9929, n_9930;
  wire n_9931, n_9932, n_9933, n_9934, n_9935, n_9936, n_9937, n_9938;
  wire n_9939, n_9940, n_9941, n_9942, n_9943, n_9944, n_9945, n_9946;
  wire n_9947, n_9948, n_9951, n_9952, n_9954, n_9955, n_9956, n_9957;
  wire n_9958, n_9959, n_9960, n_9961, n_9962, n_9963, n_9964, n_9965;
  wire n_9966, n_9967, n_9968, n_9969, n_9970, n_9971, n_9972, n_9973;
  wire n_9974, n_9975, n_9976, n_9977, n_9978, n_9979, n_9980, n_9981;
  wire n_9982, n_9983, n_9984, n_9985, n_9986, n_9987, n_9988, n_9989;
  wire n_9990, n_9991, n_9992, n_9993, n_9995, n_9996, n_9997, n_9998;
  wire n_9999, n_10000, n_10001, n_10002, n_10003, n_10004, n_10005,
       n_10006;
  wire n_10007, n_10008, n_10009, n_10010, n_10011, n_10012, n_10013,
       n_10014;
  wire n_10015, n_10016, n_10017, n_10018, n_10020, n_10021, n_10022,
       n_10023;
  wire n_10024, n_10025, n_10026, n_10027, n_10028, n_10030, n_10031,
       n_10032;
  wire n_10033, n_10034, n_10035, n_10036, n_10037, n_10038, n_10039,
       n_10040;
  wire n_10041, n_10042, n_10043, n_10044, n_10045, n_10046, n_10047,
       n_10048;
  wire n_10049, n_10050, n_10051, n_10052, n_10053, n_10054, n_10055,
       n_10056;
  wire n_10057, n_10058, n_10060, n_10061, n_10062, n_10063, n_10064,
       n_10065;
  wire n_10066, n_10068, n_10069, n_10070, n_10071, n_10072, n_10073,
       n_10074;
  wire n_10076, n_10077, n_10078, n_10079, n_10080, n_10081, n_10082,
       n_10083;
  wire n_10084, n_10085, n_10086, n_10087, n_10088, n_10089, n_10090,
       n_10091;
  wire n_10092, n_10093, n_10094, n_10095, n_10096, n_10097, n_10098,
       n_10099;
  wire n_10100, n_10101, n_10102, n_10103, n_10104, n_10105, n_10106,
       n_10107;
  wire n_10108, n_10109, n_10110, n_10111, n_10112, n_10113, n_10114,
       n_10115;
  wire n_10116, n_10118, n_10119, n_10120, n_10122, n_10123, n_10125,
       n_10126;
  wire n_10127, n_10128, n_10129, n_10130, n_10131, n_10132, n_10133,
       n_10134;
  wire n_10135, n_10136, n_10137, n_10138, n_10139, n_10140, n_10141,
       n_10142;
  wire n_10143, n_10144, n_10145, n_10146, n_10147, n_10148, n_10149,
       n_10150;
  wire n_10151, n_10152, n_10153, n_10154, n_10155, n_10156, n_10157,
       n_10158;
  wire n_10159, n_10161, n_10162, n_10163, n_10164, n_10165, n_10166,
       n_10167;
  wire n_10168, n_10169, n_10170, n_10171, n_10172, n_10173, n_10174,
       n_10175;
  wire n_10176, n_10177, n_10178, n_10179, n_10180, n_10181, n_10182,
       n_10183;
  wire n_10184, n_10185, n_10186, n_10187, n_10188, n_10189, n_10190,
       n_10191;
  wire n_10192, n_10193, n_10194, n_10195, n_10196, n_10197, n_10198,
       n_10199;
  wire n_10200, n_10201, n_10202, n_10203, n_10204, n_10205, n_10207,
       n_10208;
  wire n_10209, n_10211, n_10214, n_10217, n_10220, n_10223, n_10226,
       n_10229;
  wire n_10232, n_10235, n_10238, n_10241, n_10246, n_10247, n_10252,
       n_10253;
  wire n_10258, n_10259, n_10264, n_10265, n_10270, n_10271, n_10274,
       n_10279;
  wire n_10280, n_10283, n_10288, n_10289, n_10294, n_10295, n_10304,
       n_10305;
  wire n_10306, n_10307, n_10312, n_10313, n_10316, n_10321, n_10322,
       n_10325;
  wire n_10328, n_10333, n_10334, n_10341, n_10342, n_10343, n_10348,
       n_10349;
  wire n_10352, n_10357, n_10358, n_10367, n_10368, n_10369, n_10370,
       n_10387;
  wire n_10388, n_10389, n_10390, n_10391, n_10392, n_10393, n_10394,
       n_10397;
  wire n_10404, n_10406, n_10421, n_10422, n_10423, n_10424, n_10425,
       n_10426;
  wire n_10427, n_10434, n_10435, n_10436, n_10439, n_10450, n_10451,
       n_10452;
  wire n_10453, n_10454, n_10465, n_10466, n_10467, n_10468, n_10469,
       n_10472;
  wire n_10478, n_10481, n_10484, n_10487, n_10490, n_10493, n_10510,
       n_10511;
  wire n_10512, n_10513, n_10514, n_10515, n_10516, n_10517, n_10530,
       n_10531;
  wire n_10532, n_10533, n_10534, n_10535, n_10548, n_10549, n_10550,
       n_10551;
  wire n_10552, n_10553, n_10566, n_10567, n_10568, n_10569, n_10570,
       n_10571;
  wire n_10584, n_10585, n_10586, n_10587, n_10588, n_10589, n_10598,
       n_10599;
  wire n_10600, n_10601, n_10604, n_10607, n_10610, n_10613, n_10616,
       n_10619;
  wire n_10622, n_10625, n_10628, n_10631, n_10634, n_10637, n_10640,
       n_10647;
  wire n_10648, n_10649, n_10654, n_10655, n_10664, n_10665, n_10666,
       n_10667;
  wire n_10672, n_10673, n_10680, n_10682, n_10685, n_10692, n_10693,
       n_10694;
  wire n_10701, n_10702, n_10703, n_10706, n_10715, n_10716, n_10717,
       n_10718;
  wire n_10731, n_10732, n_10733, n_10734, n_10735, n_10736, n_10749,
       n_10750;
  wire n_10751, n_10752, n_10753, n_10754, n_10767, n_10768, n_10769,
       n_10770;
  wire n_10771, n_10772, n_10785, n_10786, n_10787, n_10788, n_10789,
       n_10790;
  wire n_10803, n_10804, n_10805, n_10806, n_10807, n_10808, n_10817,
       n_10818;
  wire n_10819, n_10820, n_10825, n_10826, n_10829, n_10832, n_10835,
       n_10838;
  wire n_10841, n_10844, n_10847, n_10850, n_10853, n_10856, n_10859,
       n_10862;
  wire n_10865, n_10868, n_10871, n_10874, n_10877, n_10880, n_10885,
       n_10886;
  wire n_10901, n_10902, n_10903, n_10904, n_10905, n_10906, n_10907,
       n_10910;
  wire n_10919, n_10920, n_10921, n_10922, n_10935, n_10936, n_10937,
       n_10938;
  wire n_10939, n_10940, n_10953, n_10954, n_10955, n_10956, n_10957,
       n_10958;
  wire n_10971, n_10972, n_10973, n_10974, n_10975, n_10976, n_10989,
       n_10990;
  wire n_10991, n_10992, n_10993, n_10994, n_11007, n_11008, n_11009,
       n_11010;
  wire n_11011, n_11012, n_11025, n_11026, n_11027, n_11028, n_11029,
       n_11030;
  wire n_11043, n_11044, n_11045, n_11046, n_11047, n_11048, n_11051,
       n_11054;
  wire n_11057, n_11060, n_11063, n_11066, n_11069, n_11072, n_11075,
       n_11078;
  wire n_11081, n_11084, n_11087, n_11090, n_11093, n_11096, n_11099,
       n_11102;
  wire n_11105, n_11108, n_11111, n_11114, n_11117, n_11124, n_11125,
       n_11126;
  wire n_11129, n_11142, n_11144, n_11149, n_11150, n_11158, n_11159,
       n_11170;
  wire n_11171, n_11172, n_11173, n_11174, n_11187, n_11188, n_11189,
       n_11190;
  wire n_11191, n_11192, n_11205, n_11206, n_11207, n_11208, n_11209,
       n_11210;
  wire n_11223, n_11224, n_11225, n_11226, n_11227, n_11228, n_11241,
       n_11242;
  wire n_11243, n_11244, n_11245, n_11246, n_11257, n_11258, n_11259,
       n_11260;
  wire n_11261, n_11274, n_11275, n_11276, n_11277, n_11278, n_11279,
       n_11292;
  wire n_11293, n_11294, n_11295, n_11296, n_11297, n_11310, n_11311,
       n_11312;
  wire n_11313, n_11314, n_11315, n_11328, n_11329, n_11330, n_11331,
       n_11332;
  wire n_11333, n_11346, n_11347, n_11348, n_11349, n_11350, n_11351,
       n_11354;
  wire n_11357, n_11360, n_11363, n_11366, n_11369, n_11372, n_11375,
       n_11378;
  wire n_11381, n_11384, n_11387, n_11390, n_11393, n_11396, n_11399,
       n_11402;
  wire n_11405, n_11408, n_11411, n_11414, n_11417, n_11420, n_11423,
       n_11426;
  wire n_11429, n_11434, n_11435, n_11438, n_11441, n_11444, n_11447,
       n_11450;
  wire n_11457, n_11458, n_11459, n_11466, n_11468, n_11483, n_11484,
       n_11485;
  wire n_11486, n_11487, n_11488, n_11489, n_11500, n_11501, n_11502,
       n_11503;
  wire n_11504, n_11509, n_11510, n_11519, n_11520, n_11521, n_11522,
       n_11535;
  wire n_11536, n_11537, n_11538, n_11539, n_11540, n_11553, n_11554,
       n_11555;
  wire n_11556, n_11557, n_11558, n_11571, n_11572, n_11573, n_11574,
       n_11575;
  wire n_11576, n_11589, n_11590, n_11591, n_11592, n_11593, n_11594,
       n_11607;
  wire n_11608, n_11609, n_11610, n_11611, n_11612, n_11625, n_11626,
       n_11627;
  wire n_11628, n_11629, n_11630, n_11643, n_11644, n_11645, n_11646,
       n_11647;
  wire n_11648, n_11661, n_11662, n_11663, n_11664, n_11665, n_11666,
       n_11679;
  wire n_11680, n_11681, n_11682, n_11683, n_11684, n_11697, n_11698,
       n_11699;
  wire n_11700, n_11701, n_11702, n_11715, n_11716, n_11717, n_11718,
       n_11719;
  wire n_11720, n_11723, n_11730, n_11731, n_11732, n_11739, n_11740,
       n_11741;
  wire n_11748, n_11749, n_11750, n_11753, n_11756, n_11763, n_11764,
       n_11765;
  wire n_11774, n_11775, n_11776, n_11777, n_11786, n_11787, n_11788,
       n_11789;
  wire n_11798, n_11799, n_11800, n_11801, n_11810, n_11811, n_11812,
       n_11813;
  wire n_11822, n_11823, n_11824, n_11825, n_11832, n_11833, n_11834,
       n_11841;
  wire n_11842, n_11843, n_11856, n_11857, n_11858, n_11859, n_11860,
       n_11861;
  wire n_11866, n_11867, n_11874, n_11875, n_11876, n_11881, n_11882,
       n_11887;
  wire n_11888, n_11895, n_11896, n_11897, n_11900, n_11905, n_11906,
       n_11915;
  wire n_11916, n_11917, n_11918, n_11925, n_11926, n_11927, n_11934,
       n_11935;
  wire n_11936, n_11947, n_11948, n_11949, n_11950, n_11951, n_11958,
       n_11959;
  wire n_11960, n_11967, n_11968, n_11969, n_11976, n_11977, n_11978,
       n_11985;
  wire n_11986, n_11987, n_11990, n_11993, n_11996, n_12001, n_12002,
       n_12009;
  wire n_12010, n_12011, n_12016, n_12017, n_12024, n_12025, n_12026,
       n_12031;
  wire n_12032, n_12037, n_12038, n_12041, n_12054, n_12055, n_12056,
       n_12057;
  wire n_12058, n_12059, n_12062, n_12069, n_12070, n_12071, n_12076,
       n_12077;
  wire n_12080, n_12085, n_12086, n_12089, n_12092, n_12095, n_12098,
       n_12101;
  wire n_12106, n_12107, n_12124, n_12125, n_12126, n_12127, n_12128,
       n_12129;
  wire n_12130, n_12131, n_12138, n_12139, n_12140, n_12143, n_12146,
       n_12149;
  wire n_12152, n_12155, n_12158, n_12161, n_12164, n_12167, n_12170,
       n_12173;
  wire n_12176, n_12179, n_12182, n_12185, n_12194, n_12195, n_12196,
       n_12197;
  wire n_12200, n_12203, n_12206, n_12209, n_12212, n_12215, n_12218,
       n_12221;
  wire n_12224, n_12227, n_12230, n_12233, n_12236, n_12239, n_12242,
       n_12245;
  wire n_12248, n_12257, n_12258, n_12259, n_12260, n_12263, n_12266,
       n_12269;
  wire n_12272, n_12275, n_12278, n_12281, n_12284, n_12287, n_12290,
       n_12293;
  wire n_12296, n_12299, n_12302, n_12305, n_12308, n_12311, n_12314,
       n_12317;
  wire n_12320, n_12323, n_12328, n_12329, n_12341, n_12342, n_12343,
       n_12344;
  wire n_12347, n_12350, n_12353, n_12356, n_12359, n_12362, n_12365,
       n_12368;
  wire n_12371, n_12374, n_12377, n_12380, n_12383, n_12386, n_12389,
       n_12392;
  wire n_12395, n_12398, n_12401, n_12404, n_12407, n_12410, n_12413,
       n_12416;
  wire n_12419, n_12422, n_12433, n_12434, n_12435, n_12436, n_12437,
       n_12634;
  wire n_12635, n_12638, n_12639, n_12640, n_12641, n_12642, n_12643,
       n_12644;
  wire n_12645, n_12646, n_12647, n_12648, n_12649, n_12650, n_12651,
       n_12652;
  wire n_12653, n_12654, n_12655, n_12656, n_12657, n_12658, n_12659,
       n_12660;
  wire n_12661, n_12662, n_12663, n_12664, n_12665, n_12666, n_12667,
       n_12668;
  wire n_12669, n_12670, n_12671, n_12672, n_12673, n_12674, n_12675,
       n_12676;
  wire n_12677, n_12678, n_12679, n_12680, n_12681, n_12682, n_12683,
       n_12684;
  wire n_12685, n_12686, n_12687, n_12688, n_12689, n_12690, n_12691,
       n_12692;
  wire n_12693, n_12694, n_12695, n_12696, n_12697, n_12698, n_12699,
       n_12700;
  wire n_12701, n_12702, n_12703, n_12706, n_12707, n_12708, n_12709,
       n_12710;
  wire n_12711, n_12712, n_12713, n_12714, n_12715, n_12716, n_12717,
       n_12718;
  wire n_12719, n_12720, n_12721, n_12722, n_12723, n_12724, n_12725,
       n_12726;
  wire n_12727, n_12728, n_12729, n_12730, n_12731, n_12732, n_12733,
       n_12734;
  wire n_12735, n_12736, n_12737, n_12738, n_12739, n_12740, n_12741,
       n_12742;
  wire n_12743, n_12744, n_12745, n_12746, n_12747, n_12748, n_12749,
       n_12750;
  wire n_12751, n_12752, n_12753, n_12754, n_12755, n_12756, n_12757,
       n_12758;
  wire n_12759, n_12762, n_12763, n_12764, n_12765, n_12766, n_12767,
       n_12768;
  wire n_12769, n_12770, n_12771, n_12772, n_12773, n_12774, n_12775,
       n_12776;
  wire n_12777, n_12778, n_12779, n_12780, n_12781, n_12782, n_12783,
       n_12784;
  wire n_12785, n_12786, n_12787, n_12788, n_12789, n_12790, n_12791,
       n_12792;
  wire n_12793, n_12794, n_12795, n_12796, n_12797, n_12798, n_12799,
       n_12800;
  wire n_12801, n_12802, n_12803, n_12804, n_12805, n_12808, n_12809,
       n_12810;
  wire n_12812, n_12813, n_12814, n_12815, n_12816, n_12817, n_12818,
       n_12819;
  wire n_12820, n_12821, n_12822, n_12823, n_12824, n_12825, n_12826,
       n_12827;
  wire n_12828, n_12829, n_12830, n_12831, n_12832, n_12833, n_12834,
       n_12835;
  wire n_12836, n_12837, n_12840, n_12842, n_12843, n_12844, n_12845,
       n_12846;
  wire n_12847, n_12848, n_12849, n_12850, n_12851, n_12852, n_12853,
       n_12854;
  wire n_12855, n_12856, n_12857, n_12860, n_12861, n_12863, n_12864,
       n_12865;
  wire n_12866, n_12867, n_12868, n_12869, n_12870, n_12871, n_12872,
       n_12873;
  wire n_12874, n_12875, n_12876, n_12877, n_12878, n_12880, n_12881,
       n_12882;
  wire n_12883, n_12884, n_12885, n_12886, n_12887, n_12888, n_12889,
       n_12890;
  wire n_12891, n_12892, n_12893, n_12894, n_12895, n_12896, n_12898,
       n_12899;
  wire n_12900, n_12901, n_12902, n_12903, n_12904, n_12905, n_12906,
       n_12907;
  wire n_12908, n_12909, n_12910, n_12911, n_12912, n_12913, n_12914,
       n_12915;
  wire n_12916, n_12917, n_12918, n_12919, n_12920, n_12921, n_12922,
       n_12923;
  wire n_12924, n_12925, n_12926, n_12927, n_12928, n_12929, n_12930,
       n_12931;
  wire n_12932, n_12933, n_12934, n_12935;
  nand anoymous (n_9353, b6, b7);
  or g16819 (n_9413, b4, wc);
  not gc (wc, n_9402);
  or g16853 (n_9429, b5, wc0);
  not gc0 (wc0, n_9428);
  or g16854 (n_9451, b6, wc1);
  not gc1 (wc1, n_9428);
  or g17045 (n_9601, b11, wc2);
  not gc2 (wc2, n_9600);
  nand g18127 (n_9730, n_9725, n_9729);
  nand g18137 (n_9709, n_9705, n_9708);
  nand g18187 (n_9359, b11, b10);
  nand g18204 (n_9347, b4, b5);
  nand g18210 (n_9343, b3, b2);
  or g18265 (n_9398, n_9397, wc3);
  not gc3 (wc3, a13);
  nand g18283 (n_9360, b12, b11);
  or g18299 (n_9320, b10, b9);
  or g18304 (n_9316, b6, b5);
  or g18306 (n_9323, n_9316, n_9322);
  or g18413 (n_9324, b1, b2);
  or g18724 (n_9339, wc4, a14);
  not gc4 (wc4, b0);
  or g18774 (n_9403, b3, wc5);
  not gc5 (wc5, n_9402);
  or g18806 (n_9430, wc6, n_9428);
  not gc6 (wc6, b5);
  or g18855 (n_9503, wc7, n_9472);
  not gc7 (wc7, b8);
  or g19092 (n_9731, wc8, n_9729);
  not gc8 (wc8, b6);
  or g22901 (n_9317, b7, b8);
  or g22902 (n_9319, b11, b12);
  or g22909 (n_9390, wc9, a12);
  not gc9 (wc9, b0);
  or g22914 (n_9414, wc10, a10);
  not gc10 (wc10, b0);
  or g22919 (n_9452, wc11, a8);
  not gc11 (wc11, b0);
  or g22926 (n_9504, wc12, a6);
  not gc12 (wc12, b0);
  or g22930 (n_9529, b9, wc13);
  not gc13 (wc13, n_9527);
  or g22931 (n_9534, b7, wc14);
  not gc14 (wc14, n_9533);
  or g22932 (n_9540, wc15, n_9533);
  not gc15 (wc15, b7);
  or g22938 (n_9572, wc16, a4);
  not gc16 (wc16, b0);
  or g22951 (n_9653, wc17, a2);
  not gc17 (wc17, b0);
  or g22955 (n_9743, wc18, a1);
  not gc18 (wc18, b0);
  or g23508 (n_9839, wc19, n_9527);
  not gc19 (wc19, n_9377);
  nand g23538 (n_9526, n_9850, n_9503);
  or g23553 (n_9856, a11, n_9414);
  nand g23565 (n_9861, n_9463, n_9469);
  or g23568 (n_9862, a3, n_9653);
  nand g23571 (n_9863, n_9677, n_9678);
  or g23574 (n_9864, a9, n_9452);
  nand g23582 (n_9867, n_9534, n_9540);
  nand g23585 (n_9868, n_9586, n_9596);
  nand g23593 (n_9871, b1, b0);
  or g23605 (n_9875, a7, n_9504);
  or g23614 (n_9879, a5, n_9572);
  or g23617 (n_9880, wc20, n_9365);
  not gc20 (wc20, n_9359);
  or g23627 (n_9884, n_9371, wc21);
  not gc21 (wc21, n_9600);
  nand g23649 (n_9894, n_9319, n_9360);
  or g23670 (n_9901, n_9743, n_9745);
  nand g23680 (n_9622, n_9904, b0);
  nand g23681 (n_9905, n_9353, n_9362);
  nand g23692 (n_9703, n_9908, n_9668);
  nand g23720 (n_9436, n_9918, b0);
  nand g23737 (n_9925, a15, n_9339);
  nand g23786 (n_9405, n_9941, b0);
  nand g23806 (n_9482, n_9948, b0);
  nand g23816 (n_9550, n_9952, b0);
  nand g23944 (n_9997, b0, n_9744);
  or g23965 (n_10000, wc22, a13);
  not gc22 (wc22, b1);
  or g23993 (n_9973, wc23, n_9409);
  not gc23 (wc23, b2);
  or g23994 (n_9972, wc24, n_9409);
  not gc24 (wc24, b3);
  or g23998 (n_9977, wc25, n_9406);
  not gc25 (wc25, b1);
  or g23999 (n_9912, wc26, n_9406);
  not gc26 (wc26, b2);
  or g24000 (n_9975, wc27, n_9406);
  not gc27 (wc27, n_9400);
  or g24021 (n_9970, wc28, n_9447);
  not gc28 (wc28, b4);
  or g24022 (n_9898, wc29, n_9434);
  not gc29 (wc29, b3);
  or g24023 (n_9951, wc30, n_9441);
  not gc30 (wc30, b2);
  or g24024 (n_9909, wc31, n_9447);
  not gc31 (wc31, b5);
  or g24025 (n_9896, wc32, n_9434);
  not gc32 (wc32, b4);
  or g24026 (n_9917, wc33, n_9441);
  not gc33 (wc33, b3);
  or g24036 (n_9920, wc34, n_9437);
  not gc34 (wc34, b1);
  or g24037 (n_9919, wc35, n_9437);
  not gc35 (wc35, b2);
  or g24038 (n_10003, wc36, n_9437);
  not gc36 (wc36, n_9400);
  or g24066 (n_9930, wc37, n_9499);
  not gc37 (wc37, b6);
  or g24067 (n_9933, wc38, n_9476);
  not gc38 (wc38, b5);
  or g24068 (n_9935, wc39, n_9493);
  not gc39 (wc39, b4);
  or g24069 (n_9939, wc40, n_9480);
  not gc40 (wc40, b3);
  or g24070 (n_9903, wc41, n_9487);
  not gc41 (wc41, b2);
  or g24071 (n_9850, b8, wc42);
  not gc42 (wc42, n_9472);
  or g24072 (n_9929, wc43, n_9499);
  not gc43 (wc43, b7);
  or g24073 (n_9906, wc44, n_9476);
  not gc44 (wc44, b6);
  or g24074 (n_9934, wc45, n_9493);
  not gc45 (wc45, b5);
  or g24075 (n_9938, wc46, n_9480);
  not gc46 (wc46, b4);
  or g24076 (n_9998, wc47, n_9487);
  not gc47 (wc47, b3);
  or g24092 (n_9984, wc48, n_9483);
  not gc48 (wc48, b1);
  or g24093 (n_9967, wc49, n_9483);
  not gc49 (wc49, b2);
  or g24094 (n_9986, wc50, n_9483);
  not gc50 (wc50, n_9400);
  or g24130 (n_9916, wc51, n_9567);
  not gc51 (wc51, b6);
  or g24131 (n_9914, wc52, n_9544);
  not gc52 (wc52, b5);
  or g24132 (n_9976, wc53, n_9561);
  not gc53 (wc53, b4);
  or g24133 (n_9960, wc54, n_9548);
  not gc54 (wc54, b3);
  or g24134 (n_9995, wc55, n_9555);
  not gc55 (wc55, b2);
  or g24135 (n_9886, wc56, n_9538);
  not gc56 (wc56, b9);
  or g24136 (n_9889, wc57, n_9533);
  not gc57 (wc57, b8);
  or g24137 (n_9946, wc58, n_9567);
  not gc58 (wc58, b7);
  or g24138 (n_9943, wc59, n_9544);
  not gc59 (wc59, b6);
  or g24139 (n_9895, wc60, n_9561);
  not gc60 (wc60, b5);
  or g24140 (n_9899, wc61, n_9548);
  not gc61 (wc61, b4);
  or g24141 (n_9924, wc62, n_9555);
  not gc62 (wc62, b3);
  or g24142 (n_9848, wc63, n_9527);
  not gc63 (wc63, b10);
  or g24162 (n_9993, wc64, n_9551);
  not gc64 (wc64, b1);
  or g24163 (n_9915, wc65, n_9551);
  not gc65 (wc65, b2);
  or g24165 (n_9955, wc66, n_9551);
  not gc66 (wc66, n_9400);
  or g24208 (n_9969, wc67, n_9648);
  not gc67 (wc67, b10);
  or g24209 (n_9980, wc68, n_9604);
  not gc68 (wc68, b9);
  or g24210 (n_10001, wc69, n_9608);
  not gc69 (wc69, b8);
  or g24211 (n_9978, wc70, n_9612);
  not gc70 (wc70, b7);
  or g24212 (n_9937, wc71, n_9639);
  not gc71 (wc71, b6);
  or g24213 (n_9999, wc72, n_9616);
  not gc72 (wc72, b5);
  or g24214 (n_9996, wc73, n_9633);
  not gc73 (wc73, b4);
  or g24215 (n_9927, wc74, n_9620);
  not gc74 (wc74, b3);
  or g24216 (n_9966, wc75, n_9627);
  not gc75 (wc75, b2);
  or g24217 (n_9841, wc76, n_9600);
  not gc76 (wc76, b12);
  or g24218 (n_9942, wc77, n_9648);
  not gc77 (wc77, b11);
  or g24219 (n_9982, wc78, n_9604);
  not gc78 (wc78, b10);
  or g24220 (n_9940, wc79, n_9608);
  not gc79 (wc79, b9);
  or g24221 (n_9990, wc80, n_9612);
  not gc80 (wc80, b8);
  or g24222 (n_9922, wc81, n_9639);
  not gc81 (wc81, b7);
  or g24223 (n_9991, wc82, n_9616);
  not gc82 (wc82, b6);
  or g24224 (n_9992, wc83, n_9633);
  not gc83 (wc83, b5);
  or g24225 (n_9928, wc84, n_9620);
  not gc84 (wc84, b4);
  or g24226 (n_9989, wc85, n_9627);
  not gc85 (wc85, b3);
  or g24252 (n_9957, wc86, n_9623);
  not gc86 (wc86, b1);
  or g24253 (n_9962, wc87, n_9623);
  not gc87 (wc87, n_9400);
  or g24254 (n_9988, wc88, n_9623);
  not gc88 (wc88, b2);
  or g24303 (n_9843, b12, wc89);
  not gc89 (wc89, n_9694);
  or g24305 (n_9852, wc90, n_9705);
  not gc90 (wc90, b10);
  or g24417 (n_9887, wc91, n_9464);
  not gc91 (wc91, n_9428);
  or g24596 (n_10005, n_9377, wc92);
  not gc92 (wc92, n_9527);
  or g24606 (n_10010, n_9352, n_9730);
  or g24614 (n_10014, n_9730, b6);
  or g24618 (n_10016, n_9700, b14);
  or g24626 (n_10020, n_9709, n_9377);
  or g24656 (n_10035, n_9739, wc93);
  not gc93 (wc93, b5);
  or g24658 (n_10036, n_9735, wc94);
  not gc94 (wc94, b4);
  or g24672 (n_10043, n_9715, wc95);
  not gc95 (wc95, b8);
  or g24674 (n_10044, n_9719, wc96);
  not gc96 (wc96, b9);
  or g24680 (n_10047, n_9698, wc97);
  not gc97 (wc97, b13);
  or g24682 (n_10048, n_9708, wc98);
  not gc98 (wc98, b9);
  or g24684 (n_10049, n_9725, wc99);
  not gc99 (wc99, b6);
  or g24686 (n_10050, n_9729, wc100);
  not gc100 (wc100, b7);
  or g24688 (n_10051, n_9705, wc101);
  not gc101 (wc101, b11);
  or g24690 (n_10052, n_9708, wc102);
  not gc102 (wc102, b10);
  or g24694 (n_10054, wc103, n_9698);
  not gc103 (wc103, n_9374);
  or g24698 (n_10056, n_9698, wc104);
  not gc104 (wc104, b14);
  nand g24706 (n_10060, n_9360, n_9694);
  or g24744 (n_10079, n_9346, wc105);
  not gc105 (wc105, n_9402);
  nand g24770 (n_10092, n_9384, b0);
  or g25539 (n_10058, n_9646, wc106);
  not gc106 (wc106, b8);
  or g25551 (n_10068, n_10069, b10);
  nand g26492 (n_10006, n_12076, n_12077);
  nand g26495 (n_12077, n_9751, n_9788);
  or g26497 (n_12071, n_12069, n_12070);
  nand g26498 (n_12070, n_9721, n_9750);
  or g26499 (n_9750, n_12059, n_9711);
  or g26500 (n_9788, n_9779, wc107);
  not gc107 (wc107, n_12041);
  nand g26501 (n_12076, n_9369, n_9774);
  or g26502 (n_9774, n_9766, wc108);
  not gc108 (wc108, n_12062);
  or g26503 (n_12059, n_12058, n_9710);
  nand g26509 (n_12057, n_12054, n_12055);
  or g26510 (n_12026, n_12025, n_9775);
  or g26511 (n_12038, wc109, n_12037);
  not gc109 (wc109, n_9773);
  or g26512 (n_12054, wc110, n_9742);
  not gc110 (wc110, n_10046);
  or g26514 (n_10046, n_12032, n_9740);
  or g26515 (n_9773, n_9772, wc111);
  not gc111 (wc111, n_12017);
  nand g26518 (n_12032, n_9749, n_12031);
  or g26519 (n_12011, n_12010, n_9782);
  or g26522 (n_12010, wc112, n_12009);
  not gc112 (wc112, n_9784);
  nand g26523 (n_9741, n_11917, n_11918);
  nand g26524 (n_9749, n_12001, n_12002);
  nand g26525 (n_11993, n_10038, n_9720);
  nand g26526 (n_9781, n_10009, n_9780);
  nand g26527 (n_9779, n_10017, n_9778);
  nand g26528 (n_9766, n_10013, n_9765);
  nand g26530 (n_9786, n_10015, n_9785);
  nand g26533 (n_9771, n_11977, n_11978);
  or g26534 (n_10011, n_11876, wc113);
  not gc113 (wc113, n_9827);
  nand g26536 (n_11960, n_9769, n_11958);
  nand g26537 (n_9761, n_11968, n_11969);
  nand g26538 (n_12016, n_10031, n_10030);
  or g26539 (n_10021, n_11897, wc114);
  not gc114 (wc114, n_9826);
  or g26540 (n_9765, wc115, n_9763);
  not gc115 (wc115, n_10025);
  nand g26541 (n_12037, n_10041, n_10040);
  or g26542 (n_9784, n_11950, n_11951);
  or g26543 (n_11918, n_11916, b3);
  or g26544 (n_10015, n_11882, wc116);
  not gc116 (wc116, n_9827);
  or g26545 (n_10034, n_11801, wc117);
  not gc117 (wc117, n_9801);
  nand g26546 (n_12002, n_10028, n_9748);
  or g26548 (n_10038, n_11825, wc118);
  not gc118 (wc118, n_9807);
  or g26550 (n_10017, n_11888, wc119);
  not gc119 (wc119, n_9822);
  or g26551 (n_9778, wc120, n_9776);
  not gc120 (wc120, n_10027);
  nand g26552 (n_12069, n_10061, n_9701);
  or g26554 (n_11969, n_11967, n_9382);
  nand g26555 (n_10025, n_11764, n_11765);
  nand g26557 (n_10041, n_9815, n_11996);
  or g26558 (n_11741, n_11740, wc121);
  not gc121 (wc121, n_9826);
  or g26559 (n_11917, n_11915, wc122);
  not gc122 (wc122, n_9739);
  or g26560 (n_10028, n_11987, wc123);
  not gc123 (wc123, b2);
  or g26562 (n_12001, wc124, b2);
  not gc124 (wc124, n_11987);
  or g26564 (n_11978, n_11976, n_9349);
  nand g26565 (n_10031, n_9812, n_11990);
  nand g26566 (n_10027, n_11905, n_11906);
  nand g26567 (n_11897, n_11895, n_11896);
  or g26569 (n_10013, n_11750, wc125);
  not gc125 (wc125, n_9822);
  nand g26571 (n_11888, n_11887, n_9851);
  or g26572 (n_11825, n_11824, wc126);
  not gc126 (wc126, n_9826);
  nand g26573 (n_11876, n_11874, n_11875);
  nand g26575 (n_11950, n_9783, n_11947);
  or g26576 (n_11801, n_11800, wc127);
  not gc127 (wc127, n_9827);
  or g26578 (n_9701, n_11732, wc128);
  not gc128 (wc128, n_9822);
  or g26579 (n_10061, n_11927, n_9699);
  nand g26580 (n_11882, n_11881, n_9731);
  or g26582 (n_9710, n_11936, n_9699);
  nand g26583 (n_11927, n_11925, n_11926);
  nand g26584 (n_11824, n_11822, n_11823);
  nand g26585 (n_11777, n_11774, n_11775);
  nand g26586 (n_11740, n_11739, n_9852);
  nand g26587 (n_11813, n_11810, n_11811);
  nand g26588 (n_11987, n_11985, n_11986);
  or g26590 (n_9777, n_11843, n_9776);
  nand g26591 (n_11800, n_11798, n_11799);
  nand g26592 (n_11915, n_10039, n_9731);
  nand g26593 (n_11905, n_10026, n_9689);
  or g26594 (n_9812, n_9346, n_9767);
  or g26595 (n_9815, n_9381, n_9760);
  nand g26596 (n_11887, n_10016, b15);
  nand g26597 (n_11750, n_11748, n_11749);
  or g26599 (n_9783, n_11860, n_11861);
  nand g26600 (n_11881, n_10014, b7);
  or g26601 (n_9764, n_11867, n_9763);
  nand g26602 (n_11895, n_10020, n_9378);
  or g26603 (n_11967, n_9760, wc129);
  not gc129 (wc129, n_9719);
  nand g26604 (n_11874, n_10010, n_9355);
  or g26605 (n_11976, n_9767, wc130);
  not gc130 (wc130, n_9739);
  or g26608 (n_11958, wc131, n_9357);
  not gc131 (wc131, n_10022);
  nand g26609 (n_11789, n_11786, n_11787);
  nand g26610 (n_11732, n_11730, n_11731);
  nand g26611 (n_9775, n_10052, n_10051);
  nand g26612 (n_11749, n_9373, n_9700);
  nand g26613 (n_11925, n_10060, n_9319);
  or g26614 (n_10022, n_9748, wc132);
  not gc132 (wc132, n_11900);
  nand g26615 (n_9776, n_10056, n_10055);
  nand g26616 (n_9760, n_10063, n_10062);
  nand g26617 (n_12436, n_12433, n_12434);
  nand g26618 (n_12009, n_10036, n_10035);
  or g26619 (n_11986, wc133, b1);
  not gc133 (wc133, n_9901);
  nand g26620 (n_11834, n_11832, n_11833);
  nand g26621 (n_11739, n_9709, b11);
  nand g26622 (n_12024, n_10044, n_10043);
  or g26623 (n_11959, n_9828, n_9400);
  nand g26624 (n_9782, n_10050, n_10049);
  nand g26625 (n_9711, n_10048, n_9852);
  nand g26626 (n_9699, n_10047, n_9851);
  nand g26627 (n_10024, n_9799, n_11756);
  nand g26628 (n_11822, n_9709, b10);
  nand g26629 (n_10026, n_9330, n_9843);
  nand g26630 (n_10039, n_9326, n_11723);
  or g26631 (n_11786, n_9799, b4);
  nand g26632 (n_11731, n_9700, b14);
  nand g26633 (n_9767, n_10065, n_10064);
  nand g26634 (n_11843, n_11841, n_11842);
  nand g26635 (n_10023, n_9792, n_11753);
  nand g26637 (n_11861, n_11858, n_11859);
  or g26638 (n_11810, n_9792, b7);
  nand g26639 (n_11936, n_11934, n_11935);
  nand g26640 (n_11867, n_11866, n_9853);
  or g26641 (n_11947, n_9828, b2);
  nand g26642 (n_9763, n_10054, n_10053);
  nand g26643 (n_11798, n_9730, b6);
  or g26644 (n_11775, n_9792, b8);
  nand g26646 (n_11951, n_11948, n_11949);
  or g26647 (n_12056, n_9715, wc134);
  not gc134 (wc134, b7);
  or g26649 (n_9700, n_9695, wc135);
  not gc135 (wc135, n_9698);
  or g26656 (n_11858, n_9748, wc136);
  not gc136 (wc136, b3);
  or g26657 (n_11859, n_9745, wc137);
  not gc137 (wc137, b2);
  or g26658 (n_11788, wc138, b5);
  not gc138 (wc138, n_9739);
  or g26662 (n_11833, n_9725, wc139);
  not gc139 (wc139, b5);
  or g26664 (n_11811, n_9317, wc140);
  not gc140 (wc140, n_9715);
  nand g26665 (n_9792, n_9715, n_9719);
  or g26666 (n_11812, wc141, b8);
  not gc141 (wc141, n_9719);
  or g26667 (n_11935, n_9694, wc142);
  not gc142 (wc142, b12);
  or g26668 (n_12031, n_9735, wc143);
  not gc143 (wc143, b3);
  or g26669 (n_9826, n_9705, n_9708);
  or g26670 (n_11823, n_9705, wc144);
  not gc144 (wc144, b9);
  nand g26671 (n_9828, n_9745, n_9748);
  nand g26672 (n_9799, n_9735, n_9739);
  or g26673 (n_11934, n_9689, wc145);
  not gc145 (wc145, b11);
  or g26675 (n_11949, wc146, b3);
  not gc146 (wc146, n_9748);
  or g26676 (n_12055, n_9719, wc147);
  not gc147 (wc147, b8);
  or g26677 (n_11841, n_9689, wc148);
  not gc148 (wc148, b12);
  or g26678 (n_11842, n_9694, wc149);
  not gc149 (wc149, b13);
  or g26679 (n_11723, wc150, b4);
  not gc150 (wc150, n_9725);
  or g26680 (n_9827, n_9725, n_9729);
  or g26681 (n_11906, wc151, b13);
  not gc151 (wc151, n_9694);
  or g26682 (n_11799, n_9729, wc152);
  not gc152 (wc152, b5);
  nand g26683 (n_11985, n_9743, n_9745);
  or g26684 (n_11832, n_9739, wc153);
  not gc153 (wc153, b4);
  or g26685 (n_9822, wc154, n_9698);
  not gc154 (wc154, n_9695);
  or g26686 (n_11776, wc155, b9);
  not gc155 (wc155, n_9719);
  or g26687 (n_9748, n_11557, n_11558);
  nand g26688 (n_12634, n_9997, a2);
  or g26689 (n_12635, n_9997, a2);
  nand g26690 (n_9745, n_12634, n_12635);
  or g26691 (n_9715, n_11611, n_11612);
  or g26692 (n_9735, n_11701, n_11702);
  or g26694 (n_9719, n_11683, n_11684);
  or g26695 (n_9739, n_11719, n_11720);
  or g26696 (n_9694, n_11665, n_11666);
  or g26697 (n_9689, n_11575, n_11576);
  or g26698 (n_9725, n_11593, n_11594);
  or g26699 (n_9708, n_11539, n_11540);
  or g26700 (n_9729, n_11629, n_11630);
  or g26701 (n_9705, n_11647, n_11648);
  nand g26702 (n_11665, n_11661, n_11662);
  nand g26703 (n_11522, n_11519, n_11520);
  nand g26704 (n_11575, n_11571, n_11572);
  nand g26707 (n_11539, n_11535, n_11536);
  nand g26708 (n_11683, n_11679, n_11680);
  nand g26709 (n_11748, n_10012, n_9374);
  nand g26710 (n_11557, n_11553, n_11554);
  nand g26711 (n_11611, n_11607, n_11608);
  nand g26712 (n_11701, n_11697, n_11698);
  nand g26713 (n_11647, n_11643, n_11644);
  nand g26714 (n_11730, n_10008, b13);
  nand g26715 (n_11593, n_11589, n_11590);
  nand g26716 (n_11629, n_11625, n_11626);
  nand g26717 (n_11719, n_11715, n_11716);
  nand g26719 (n_11666, n_11663, n_11664);
  nand g26722 (n_9851, n_9695, b14);
  nand g26723 (n_10055, n_9695, b15);
  nand g26724 (n_11648, n_11645, n_11646);
  nand g26725 (n_11630, n_11627, n_11628);
  nand g26726 (n_9744, n_9666, n_9687);
  nand g26727 (n_11720, n_11717, n_11718);
  nand g26731 (n_11540, n_11537, n_11538);
  or g26732 (n_10012, n_9373, n_9695);
  nand g26734 (n_11558, n_11555, n_11556);
  nand g26735 (n_11612, n_11609, n_11610);
  nand g26736 (n_11594, n_11591, n_11592);
  nand g26737 (n_11684, n_11681, n_11682);
  nand g26741 (n_10053, n_9373, n_9695);
  nand g26742 (n_11576, n_11573, n_11574);
  nand g26745 (n_11702, n_11699, n_11700);
  or g26746 (n_10008, n_9695, b14);
  nand g26747 (n_11700, n_9623, n_9665);
  nand g26748 (n_11664, n_9648, n_9665);
  nand g26749 (n_11521, n_9600, n_9665);
  nand g26750 (n_11556, n_9665, a3);
  nand g26751 (n_11538, n_9612, n_9665);
  or g26752 (n_9666, n_9665, wc156);
  not gc156 (wc156, n_9650);
  nand g26753 (n_11592, n_9620, n_9665);
  nand g26755 (n_11610, n_9616, n_9665);
  nand g26756 (n_11646, n_9608, n_9665);
  nand g26757 (n_11574, n_9604, n_9665);
  nand g26758 (n_11718, n_9627, n_9665);
  nand g26759 (n_11682, n_9639, n_9665);
  nand g26760 (n_11628, n_9633, n_9665);
  or g26761 (n_11609, wc157, n_9688);
  not gc157 (wc157, n_10095);
  or g26762 (n_11699, wc158, n_9688);
  not gc158 (wc158, n_10110);
  or g26763 (n_11681, wc159, n_9688);
  not gc159 (wc159, n_10107);
  or g26764 (n_11717, wc160, n_9688);
  not gc160 (wc160, n_10113);
  or g26765 (n_11645, wc161, n_9688);
  not gc161 (wc161, n_10101);
  or g26766 (n_11573, wc162, n_9688);
  not gc162 (wc162, n_10086);
  or g26767 (n_11591, wc163, n_9688);
  not gc163 (wc163, n_10089);
  or g26768 (n_9665, wc164, n_9331);
  not gc164 (wc164, n_10211);
  or g26769 (n_11555, wc165, n_9688);
  not gc165 (wc165, n_10083);
  or g26770 (n_11663, wc166, n_9688);
  not gc166 (wc166, n_10104);
  or g26771 (n_11537, wc167, n_9688);
  not gc167 (wc167, n_10080);
  or g26772 (n_11627, wc168, n_9688);
  not gc168 (wc168, n_10098);
  or g26773 (n_11520, wc169, n_9688);
  not gc169 (wc169, n_10076);
  nand g26776 (n_10211, n_11509, n_11510);
  or g26789 (n_11510, wc170, n_9583);
  not gc170 (wc170, n_10209);
  or g26790 (n_9650, n_11489, b15);
  or g26791 (n_9687, n_11504, n_9373);
  or g26792 (n_11489, n_11488, n_9318);
  or g26793 (n_10209, n_11468, wc171);
  not gc171 (wc171, b13);
  or g26794 (n_11504, n_11503, wc172);
  not gc172 (wc172, n_9369);
  or g26795 (n_11509, wc173, b13);
  not gc173 (wc173, n_11468);
  or g26796 (n_11488, wc174, n_11487);
  not gc174 (wc174, n_11486);
  or g26797 (n_11503, n_11502, n_9374);
  nand g26798 (n_11468, n_11466, n_11384);
  nand g26799 (n_11502, n_11500, n_11501);
  nand g26800 (n_11466, n_9841, n_9664);
  nand g26801 (n_12638, n_9697, n_9664);
  or g26802 (n_12639, n_9697, n_9664);
  nand g26803 (n_10077, n_12638, n_12639);
  nand g26804 (n_12640, n_9696, n_9649);
  or g26805 (n_12641, n_9696, n_9649);
  nand g26806 (n_10076, n_12640, n_12641);
  or g26807 (n_11486, n_11483, n_9649);
  nand g26808 (n_9664, n_11408, n_12395);
  nand g26809 (n_9649, n_11405, n_12392);
  nand g26810 (n_11500, n_10208, n_9831);
  nand g26811 (n_12642, n_9690, n_9643);
  or g26812 (n_12643, n_9690, n_9643);
  nand g26813 (n_10104, n_12642, n_12643);
  nand g26814 (n_12392, n_9969, n_9643);
  nand g26815 (n_12395, n_9942, n_9663);
  nand g26816 (n_10208, n_11458, n_11459);
  nand g26817 (n_12644, n_9691, n_9663);
  or g26818 (n_12645, n_9691, n_9663);
  nand g26819 (n_10106, n_12644, n_12645);
  nand g26821 (n_12646, n_9693, n_9692);
  or g26822 (n_12647, n_9693, n_9692);
  nand g26823 (n_10105, n_12646, n_12647);
  nand g26824 (n_9643, n_11402, n_12389);
  nand g26825 (n_9663, n_11399, n_12386);
  nand g26826 (n_12389, n_9980, n_9642);
  nand g26827 (n_12386, n_9982, n_9662);
  or g26828 (n_9693, n_11450, wc175);
  not gc175 (wc175, n_9667);
  nand g26829 (n_12648, n_9682, n_9642);
  or g26830 (n_12649, n_9682, n_9642);
  nand g26831 (n_10086, n_12648, n_12649);
  nand g26832 (n_12650, n_9681, n_9662);
  or g26833 (n_12651, n_9681, n_9662);
  nand g26834 (n_10088, n_12650, n_12651);
  nand g26835 (n_11457, n_9685, n_9884);
  nand g26836 (n_9642, n_11387, n_12374);
  nand g26837 (n_12652, n_9680, n_9874);
  or g26838 (n_12653, n_9680, n_9874);
  nand g26839 (n_10087, n_12652, n_12653);
  nand g26840 (n_11450, n_9838, n_9684);
  or g26841 (n_9685, wc176, n_9684);
  not gc176 (wc176, n_9683);
  nand g26842 (n_9662, n_11390, n_12377);
  nand g26843 (n_12654, n_9702, n_9641);
  or g26844 (n_12655, n_9702, n_9641);
  nand g26845 (n_10101, n_12654, n_12655);
  nand g26847 (n_12656, n_9863, n_9703);
  or g26848 (n_12657, n_9863, n_9703);
  nand g26849 (n_10102, n_12656, n_12657);
  nand g26850 (n_9680, n_9679, n_11447);
  nand g26851 (n_12377, n_9940, n_9661);
  nand g26852 (n_12658, n_9704, n_9661);
  or g26853 (n_12659, n_9704, n_9661);
  nand g26854 (n_10103, n_12658, n_12659);
  nand g26855 (n_12374, n_10001, n_9641);
  nand g26856 (n_9641, n_11396, n_12383);
  nand g26858 (n_9661, n_11393, n_12380);
  nand g26859 (n_12660, n_9873, n_9676);
  or g26860 (n_12661, n_9873, n_9676);
  nand g26861 (n_10081, n_12660, n_12661);
  nand g26862 (n_12662, n_9706, n_9660);
  or g26863 (n_12663, n_9706, n_9660);
  nand g26864 (n_10082, n_12662, n_12663);
  nand g26865 (n_12664, n_9707, n_9640);
  or g26866 (n_12665, n_9707, n_9640);
  nand g26867 (n_10080, n_12664, n_12665);
  nand g26868 (n_12383, n_9978, n_9640);
  nand g26869 (n_12380, n_9990, n_9660);
  nand g26870 (n_9677, n_9669, n_9676);
  nand g26871 (n_9676, n_11360, n_12350);
  nand g26872 (n_9640, n_11417, n_12404);
  nand g26873 (n_9660, n_11420, n_12407);
  nand g26874 (n_12666, n_9717, n_9675);
  or g26875 (n_12667, n_9717, n_9675);
  nand g26876 (n_10108, n_12666, n_12667);
  nand g26877 (n_12407, n_9922, n_9659);
  nand g26878 (n_12668, n_9716, n_9635);
  or g26879 (n_12669, n_9716, n_9635);
  nand g26880 (n_10107, n_12668, n_12669);
  nand g26881 (n_12404, n_9937, n_9635);
  nand g26882 (n_12670, n_9718, n_9659);
  or g26883 (n_12671, n_9718, n_9659);
  nand g26884 (n_10109, n_12670, n_12671);
  nand g26885 (n_12350, n_9983, n_9675);
  nand g26886 (n_9675, n_11363, n_12353);
  nand g26887 (n_9635, n_11414, n_12401);
  nand g26888 (n_9659, n_11411, n_12398);
  nand g26889 (n_12353, n_9979, n_9674);
  nand g26890 (n_12672, n_9714, n_9674);
  or g26891 (n_12673, n_9714, n_9674);
  nand g26892 (n_10096, n_12672, n_12673);
  nand g26893 (n_12398, n_9991, n_9658);
  nand g26894 (n_12674, n_9712, n_9658);
  or g26895 (n_12675, n_9712, n_9658);
  nand g26896 (n_10097, n_12674, n_12675);
  nand g26897 (n_12401, n_9999, n_9634);
  nand g26898 (n_12676, n_9713, n_9634);
  or g26899 (n_12677, n_9713, n_9634);
  nand g26900 (n_10095, n_12676, n_12677);
  nand g26901 (n_9674, n_11366, n_12356);
  nand g26902 (n_9634, n_11423, n_12410);
  nand g26903 (n_9658, n_11426, n_12413);
  nand g26904 (n_12356, n_9985, n_9673);
  nand g26905 (n_12678, n_9727, n_9673);
  or g26906 (n_12679, n_9727, n_9673);
  nand g26907 (n_10099, n_12678, n_12679);
  nand g26908 (n_12680, n_9657, n_9728);
  or g26909 (n_12681, n_9657, n_9728);
  nand g26910 (n_10100, n_12680, n_12681);
  nand g26911 (n_12413, n_9992, n_9657);
  nand g26912 (n_12410, n_9996, n_9629);
  nand g26913 (n_12682, n_9629, n_9726);
  or g26914 (n_12683, n_9629, n_9726);
  nand g26915 (n_10098, n_12682, n_12683);
  nand g26916 (n_9673, n_11369, n_12359);
  nand g26917 (n_9686, n_9683, n_11435);
  nand g26918 (n_9629, n_11372, n_12362);
  nand g26919 (n_9657, n_11375, n_12365);
  nand g26920 (n_12365, n_9928, n_9656);
  nand g26921 (n_12684, n_9724, n_9656);
  or g26922 (n_12685, n_9724, n_9656);
  nand g26923 (n_10091, n_12684, n_12685);
  or g26924 (n_11435, n_11434, wc177);
  not gc177 (wc177, n_9667);
  nand g26925 (n_12686, n_9723, n_9628);
  or g26926 (n_12687, n_9723, n_9628);
  nand g26927 (n_10089, n_12686, n_12687);
  nand g26928 (n_12362, n_9927, n_9628);
  nand g26929 (n_12688, n_9722, n_9672);
  or g26930 (n_12689, n_9722, n_9672);
  nand g26931 (n_10090, n_12688, n_12689);
  nand g26932 (n_12359, n_9902, n_9672);
  nand g26933 (n_9656, n_11381, n_12371);
  nand g26934 (n_11434, n_9838, n_9881);
  nand g26935 (n_9672, n_11357, n_12347);
  nand g26936 (n_9628, n_11378, n_12368);
  nand g26938 (n_12690, n_9737, n_9671);
  or g26939 (n_12691, n_9737, n_9671);
  nand g26940 (n_10114, n_12690, n_12691);
  nand g26941 (n_12368, n_9966, n_9624);
  nand g26942 (n_12347, n_9964, n_9671);
  nand g26943 (n_12692, n_9738, n_9655);
  or g26944 (n_12693, n_9738, n_9655);
  nand g26945 (n_10115, n_12692, n_12693);
  nand g26946 (n_11487, n_11484, n_11485);
  nand g26947 (n_12371, n_9989, n_9655);
  nand g26948 (n_12694, n_9736, n_9624);
  or g26949 (n_12695, n_9736, n_9624);
  nand g26950 (n_10113, n_12694, n_12695);
  nand g26951 (n_9655, n_11444, n_12422);
  nand g26952 (n_12696, n_9654, n_9734);
  or g26953 (n_12697, n_9654, n_9734);
  nand g26954 (n_10112, n_12696, n_12697);
  nand g26955 (n_9671, n_11438, n_12416);
  or g26956 (n_12698, n_9621, n_9733);
  nand g26957 (n_12699, n_9621, n_9733);
  nand g26958 (n_10110, n_12698, n_12699);
  nand g26959 (n_12700, n_9670, n_9732);
  or g26960 (n_12701, n_9670, n_9732);
  nand g26961 (n_10111, n_12700, n_12701);
  nand g26962 (n_9679, n_9668, n_11429);
  nand g26963 (n_9624, n_11441, n_12419);
  nand g26964 (n_11484, n_10071, n_9583);
  nand g26965 (n_12419, n_9621, n_9957);
  nand g26966 (n_9722, n_9902, n_11369);
  nand g26968 (n_9691, n_9942, n_11408);
  nand g26969 (n_11483, n_9958, n_9601);
  nand g26970 (n_9681, n_9982, n_11399);
  nand g26971 (n_9713, n_9999, n_11414);
  nand g26972 (n_9874, n_9652, n_9667);
  nand g26973 (n_9714, n_9979, n_11363);
  nand g26974 (n_9712, n_9991, n_11411);
  nand g26975 (n_9692, n_9683, n_9881);
  nand g26976 (n_9724, n_9928, n_11375);
  nand g26977 (n_9734, n_9988, n_11444);
  nand g26978 (n_12416, n_9670, n_9962);
  nand g26979 (n_12422, n_9654, n_9988);
  nand g26980 (n_9682, n_9980, n_11402);
  nand g26981 (n_9690, n_9969, n_11405);
  nand g26982 (n_9736, n_9966, n_11378);
  nand g26983 (n_9737, n_9964, n_11357);
  nand g26984 (n_9716, n_9937, n_11417);
  nand g26985 (n_9717, n_9983, n_11360);
  nand g26986 (n_9718, n_9922, n_11420);
  nand g26987 (n_9707, n_9978, n_11396);
  or g26988 (n_11485, n_9841, wc178);
  not gc178 (wc178, b11);
  nand g26989 (n_9697, n_9841, n_11384);
  nand g26990 (n_9873, n_9669, n_9678);
  nand g26991 (n_9696, n_11354, n_9601);
  nand g26992 (n_9706, n_9990, n_11393);
  nand g26993 (n_9738, n_9989, n_11381);
  nand g26994 (n_9733, n_9957, n_11441);
  nand g26995 (n_11429, n_9678, n_9908);
  nand g26996 (n_9702, n_10001, n_11387);
  nand g26997 (n_9704, n_9940, n_11390);
  nand g26998 (n_9726, n_9996, n_11423);
  nand g26999 (n_9723, n_9927, n_11372);
  nand g27000 (n_9728, n_9992, n_11426);
  nand g27001 (n_9732, n_9962, n_11438);
  nand g27002 (n_9727, n_9985, n_11366);
  or g27004 (n_11384, wc179, b12);
  not gc179 (wc179, n_9600);
  or g27005 (n_11417, wc180, b6);
  not gc180 (wc180, n_9639);
  or g27006 (n_11396, wc181, b7);
  not gc181 (wc181, n_9612);
  or g27007 (n_11387, wc182, b8);
  not gc182 (wc182, n_9608);
  or g27014 (n_11438, wc183, n_9400);
  not gc183 (wc183, n_9623);
  or g27015 (n_11378, wc184, b2);
  not gc184 (wc184, n_9627);
  or g27016 (n_11441, wc185, b1);
  not gc185 (wc185, n_9623);
  or g27017 (n_11444, wc186, b2);
  not gc186 (wc186, n_9623);
  or g27018 (n_11381, wc187, b3);
  not gc187 (wc187, n_9627);
  or g27019 (n_11375, wc188, b4);
  not gc188 (wc188, n_9620);
  or g27020 (n_11426, wc189, b5);
  not gc189 (wc189, n_9633);
  or g27021 (n_11411, wc190, b6);
  not gc190 (wc190, n_9616);
  or g27022 (n_11420, wc191, b7);
  not gc191 (wc191, n_9639);
  or g27023 (n_11393, wc192, b8);
  not gc192 (wc192, n_9612);
  or g27024 (n_11390, wc193, b9);
  not gc193 (wc193, n_9608);
  or g27025 (n_11399, wc194, b10);
  not gc194 (wc194, n_9604);
  or g27027 (n_11408, wc195, b11);
  not gc195 (wc195, n_9648);
  or g27028 (n_11402, wc196, b9);
  not gc196 (wc196, n_9604);
  or g27029 (n_11458, wc197, n_9600);
  not gc197 (wc197, n_9371);
  or g27030 (n_11372, wc198, b3);
  not gc198 (wc198, n_9620);
  or g27031 (n_11414, wc199, b5);
  not gc199 (wc199, n_9616);
  or g27032 (n_11354, n_9600, wc200);
  not gc200 (wc200, b11);
  or g27033 (n_11405, wc201, b10);
  not gc201 (wc201, n_9648);
  or g27034 (n_11423, wc202, b4);
  not gc202 (wc202, n_9633);
  nand g27035 (n_12702, n_9622, a4);
  or g27036 (n_12703, n_9622, a4);
  nand g27037 (n_9623, n_12702, n_12703);
  or g27038 (n_9627, n_11278, n_11279);
  or g27039 (n_9620, n_11332, n_11333);
  or g27040 (n_9633, n_11314, n_11315);
  or g27041 (n_9616, n_11296, n_11297);
  or g27042 (n_9639, n_11350, n_11351);
  or g27043 (n_9612, n_11245, n_11246);
  or g27044 (n_9608, n_11227, n_11228);
  or g27045 (n_9604, n_11209, n_11210);
  or g27046 (n_9648, n_11191, n_11192);
  nand g27048 (n_11315, n_11312, n_11313);
  nand g27049 (n_11228, n_11225, n_11226);
  nand g27050 (n_11351, n_11348, n_11349);
  nand g27051 (n_11333, n_11330, n_11331);
  nand g27052 (n_11191, n_11187, n_11188);
  nand g27053 (n_11209, n_11205, n_11206);
  nand g27054 (n_11314, n_11310, n_11311);
  nand g27055 (n_11296, n_11292, n_11293);
  nand g27056 (n_11279, n_11276, n_11277);
  nand g27057 (n_11332, n_11328, n_11329);
  nand g27058 (n_11210, n_11207, n_11208);
  nand g27059 (n_11246, n_11243, n_11244);
  nand g27060 (n_11350, n_11346, n_11347);
  nand g27061 (n_11278, n_11274, n_11275);
  nand g27062 (n_11261, n_11258, n_11259);
  nand g27063 (n_11192, n_11189, n_11190);
  nand g27066 (n_11227, n_11223, n_11224);
  nand g27067 (n_11245, n_11241, n_11242);
  nand g27068 (n_11297, n_11294, n_11295);
  or g27069 (n_11241, wc203, n_9584);
  not gc203 (wc203, n_10143);
  or g27070 (n_11310, wc204, n_9584);
  not gc204 (wc204, n_10173);
  or g27071 (n_11207, wc205, n_9598);
  not gc205 (wc205, n_10129);
  or g27072 (n_11328, wc206, n_9584);
  not gc206 (wc206, n_10176);
  or g27073 (n_11225, wc207, n_9598);
  not gc207 (wc207, n_10135);
  or g27074 (n_11294, wc208, n_9598);
  not gc208 (wc208, n_10165);
  or g27075 (n_11312, wc209, n_9598);
  not gc209 (wc209, n_10171);
  or g27076 (n_11243, wc210, n_9598);
  not gc210 (wc210, n_10141);
  nand g27077 (n_9904, n_9584, n_9597);
  or g27078 (n_11330, wc211, n_9598);
  not gc211 (wc211, n_10174);
  or g27079 (n_11260, n_11257, n_9598);
  or g27080 (n_11223, wc212, n_9584);
  not gc212 (wc212, n_10137);
  or g27081 (n_11292, wc213, n_9584);
  not gc213 (wc213, n_10167);
  or g27082 (n_11276, wc214, n_9598);
  not gc214 (wc214, n_10150);
  or g27083 (n_11258, wc215, n_9584);
  not gc215 (wc215, n_10122);
  or g27084 (n_11348, wc216, n_9598);
  not gc216 (wc216, n_10198);
  or g27085 (n_11187, wc217, n_9584);
  not gc217 (wc217, n_10128);
  or g27086 (n_11189, wc218, n_9598);
  not gc218 (wc218, n_10126);
  or g27087 (n_11346, wc219, n_9584);
  not gc219 (wc219, n_10200);
  or g27088 (n_11274, wc220, n_9584);
  not gc220 (wc220, n_10152);
  or g27089 (n_11205, wc221, n_9584);
  not gc221 (wc221, n_10131);
  or g27094 (n_9570, n_11174, b15);
  or g27095 (n_11174, n_11173, n_9319);
  or g27096 (n_9958, n_9583, b12);
  nand g27097 (n_11501, n_9583, n_9372);
  or g27098 (n_9831, n_9583, n_9372);
  or g27099 (n_11173, n_11172, n_9318);
  nand g27100 (n_11226, n_9567, n_9582);
  nand g27101 (n_11331, n_9551, n_9582);
  nand g27102 (n_11244, n_9544, n_9582);
  nand g27103 (n_11208, n_9533, n_9582);
  nand g27104 (n_11190, n_9538, n_9582);
  nand g27105 (n_11349, n_9561, n_9582);
  nand g27106 (n_11259, n_9527, n_9582);
  nand g27107 (n_11313, n_9555, n_9582);
  nand g27108 (n_11277, n_9582, a5);
  nand g27110 (n_11295, n_9548, n_9582);
  nand g27111 (n_11172, n_11170, n_11171);
  nand g27112 (n_11171, n_10068, n_9513);
  or g27113 (n_9582, wc222, n_9332);
  not gc222 (wc222, n_10207);
  nand g27114 (n_10207, n_11158, n_11159);
  nand g27115 (n_11170, n_10069, b10);
  nand g27116 (n_10069, n_9528, n_9818);
  or g27125 (n_11159, wc223, n_9513);
  not gc223 (wc223, n_10205);
  or g27127 (n_11158, wc224, b11);
  not gc224 (wc224, n_11144);
  or g27128 (n_10205, n_11144, wc225);
  not gc225 (wc225, b11);
  or g27129 (n_9597, n_11150, wc226);
  not gc226 (wc226, n_9369);
  or g27130 (n_11257, n_9529, wc227);
  not gc227 (wc227, n_9866);
  or g27131 (n_9818, wc228, n_9866);
  not gc228 (wc228, n_9529);
  nand g27132 (n_11144, n_11142, n_11072);
  or g27133 (n_11150, wc229, n_9375);
  not gc229 (wc229, n_11149);
  nand g27135 (n_11149, n_10204, n_9588);
  nand g27136 (n_11142, n_9848, n_9581);
  nand g27137 (n_12344, n_12341, n_12342);
  nand g27138 (n_12706, n_9599, n_9581);
  or g27139 (n_12707, n_9599, n_9581);
  nand g27140 (n_10122, n_12706, n_12707);
  nand g27141 (n_9581, n_11075, n_12281);
  nand g27142 (n_12342, n_10058, n_9538);
  nand g27144 (n_12281, n_9886, n_9580);
  nand g27145 (n_12708, n_9647, n_9580);
  or g27146 (n_12709, n_9647, n_9580);
  nand g27147 (n_10128, n_12708, n_12709);
  nand g27148 (n_12710, n_9644, n_9646);
  or g27149 (n_12711, n_9644, n_9646);
  nand g27150 (n_10126, n_12710, n_12711);
  nand g27152 (n_12712, n_9645, n_9868);
  or g27153 (n_12713, n_9645, n_9868);
  nand g27154 (n_10127, n_12712, n_12713);
  nand g27156 (n_9646, n_9534, n_11129);
  or g27157 (n_12341, n_11129, b8);
  nand g27158 (n_9580, n_11078, n_12284);
  nand g27159 (n_12714, n_9603, n_9579);
  or g27160 (n_12715, n_9603, n_9579);
  nand g27161 (n_10131, n_12714, n_12715);
  nand g27162 (n_9596, n_11060, n_9595);
  nand g27163 (n_12716, n_9602, n_9595);
  or g27164 (n_12717, n_9602, n_9595);
  nand g27165 (n_10130, n_12716, n_12717);
  nand g27166 (n_11129, n_9540, n_9568);
  nand g27167 (n_12718, n_9867, n_9568);
  or g27168 (n_12719, n_9867, n_9568);
  nand g27169 (n_10129, n_12718, n_12719);
  nand g27170 (n_12284, n_9889, n_9579);
  nand g27171 (n_9579, n_11081, n_12287);
  nand g27172 (n_9595, n_11057, n_12269);
  nand g27173 (n_9568, n_11084, n_12290);
  nand g27174 (n_12720, n_9605, n_9578);
  or g27175 (n_12721, n_9605, n_9578);
  nand g27176 (n_10137, n_12720, n_12721);
  nand g27177 (n_12290, n_9916, n_9563);
  nand g27178 (n_12269, n_9954, n_9594);
  nand g27179 (n_12722, n_9606, n_9594);
  or g27180 (n_12723, n_9606, n_9594);
  nand g27181 (n_10136, n_12722, n_12723);
  nand g27182 (n_12724, n_9607, n_9563);
  or g27183 (n_12725, n_9607, n_9563);
  nand g27184 (n_10135, n_12724, n_12725);
  nand g27185 (n_12287, n_9946, n_9578);
  nand g27186 (n_9594, n_11063, n_12272);
  nand g27187 (n_9563, n_11090, n_12296);
  nand g27188 (n_9578, n_11087, n_12293);
  nand g27189 (n_12726, n_9609, n_9577);
  or g27190 (n_12727, n_9609, n_9577);
  nand g27191 (n_10143, n_12726, n_12727);
  nand g27192 (n_12728, n_9611, n_9593);
  or g27193 (n_12729, n_9611, n_9593);
  nand g27194 (n_10142, n_12728, n_12729);
  nand g27195 (n_12730, n_9610, n_9562);
  or g27196 (n_12731, n_9610, n_9562);
  nand g27197 (n_10141, n_12730, n_12731);
  nand g27198 (n_12272, n_9910, n_9593);
  nand g27199 (n_12296, n_9914, n_9562);
  nand g27200 (n_12293, n_9943, n_9577);
  nand g27201 (n_9593, n_11054, n_12266);
  nand g27202 (n_9577, n_11093, n_12299);
  nand g27203 (n_9562, n_11096, n_12302);
  nand g27204 (n_12732, n_9638, n_9557);
  or g27205 (n_12733, n_9638, n_9557);
  nand g27206 (n_10198, n_12732, n_12733);
  nand g27207 (n_12266, n_9897, n_9592);
  nand g27208 (n_12734, n_9636, n_9592);
  or g27209 (n_12735, n_9636, n_9592);
  nand g27210 (n_10199, n_12734, n_12735);
  nand g27211 (n_12299, n_9895, n_9576);
  nand g27212 (n_12736, n_9637, n_9576);
  or g27213 (n_12737, n_9637, n_9576);
  nand g27214 (n_10200, n_12736, n_12737);
  nand g27215 (n_12302, n_9976, n_9557);
  nand g27216 (n_9557, n_11102, n_12308);
  nand g27217 (n_9592, n_11066, n_12275);
  nand g27218 (n_9576, n_11099, n_12305);
  nand g27219 (n_12738, n_9614, n_9556);
  or g27220 (n_12739, n_9614, n_9556);
  nand g27221 (n_10165, n_12738, n_12739);
  nand g27222 (n_9588, n_11125, n_11126);
  nand g27223 (n_12275, n_9907, n_9591);
  nand g27224 (n_12740, n_9615, n_9591);
  or g27225 (n_12741, n_9615, n_9591);
  nand g27226 (n_10166, n_12740, n_12741);
  nand g27227 (n_12305, n_9899, n_9575);
  nand g27228 (n_12742, n_9613, n_9575);
  or g27229 (n_12743, n_9613, n_9575);
  nand g27230 (n_10167, n_12742, n_12743);
  nand g27231 (n_12308, n_9960, n_9556);
  or g27232 (n_11126, wc230, n_11124);
  not gc230 (wc230, n_9587);
  nand g27233 (n_9556, n_11105, n_12311);
  nand g27234 (n_9575, n_11108, n_12314);
  nand g27235 (n_9591, n_11069, n_12278);
  nand g27236 (n_12744, n_9552, n_9630);
  or g27237 (n_12745, n_9552, n_9630);
  nand g27238 (n_10171, n_12744, n_12745);
  nand g27239 (n_12278, n_9961, n_9590);
  nand g27240 (n_12746, n_9631, n_9590);
  or g27241 (n_12747, n_9631, n_9590);
  nand g27242 (n_10172, n_12746, n_12747);
  nand g27243 (n_12748, n_9574, n_9632);
  or g27244 (n_12749, n_9574, n_9632);
  nand g27245 (n_10173, n_12748, n_12749);
  nand g27246 (n_12314, n_9924, n_9574);
  nand g27247 (n_12311, n_9995, n_9552);
  nand g27248 (n_9587, n_10007, n_9839);
  nand g27249 (n_12750, n_9589, n_9619);
  or g27250 (n_12751, n_9589, n_9619);
  nand g27251 (n_10175, n_12750, n_12751);
  nand g27252 (n_10007, n_11051, n_12263);
  nand g27253 (n_9574, n_11111, n_12317);
  nand g27254 (n_12752, n_9573, n_9617);
  or g27255 (n_12753, n_9573, n_9617);
  nand g27256 (n_10176, n_12752, n_12753);
  nand g27257 (n_9590, n_11117, n_12323);
  or g27258 (n_12754, n_9549, n_9618);
  nand g27259 (n_12755, n_9549, n_9618);
  nand g27260 (n_10174, n_12754, n_12755);
  nand g27261 (n_9552, n_11114, n_12320);
  nand g27262 (n_9615, n_9907, n_11066);
  nand g27263 (n_9605, n_9946, n_11081);
  nand g27264 (n_9618, n_9993, n_11114);
  nand g27265 (n_9613, n_9899, n_11099);
  nand g27266 (n_9599, n_9848, n_11072);
  nand g27267 (n_12323, n_9589, n_9955);
  nand g27268 (n_9606, n_9954, n_11057);
  nand g27269 (n_12320, n_9549, n_9993);
  nand g27270 (n_9614, n_9960, n_11102);
  nand g27271 (n_9630, n_9995, n_11105);
  or g27272 (n_12263, wc231, n_9586);
  not gc231 (wc231, n_9585);
  nand g27273 (n_9638, n_9976, n_11096);
  nand g27274 (n_9636, n_9897, n_11054);
  nand g27275 (n_9607, n_9916, n_11084);
  nand g27276 (n_9637, n_9895, n_11093);
  nand g27277 (n_9602, n_9586, n_11060);
  nand g27278 (n_9609, n_9943, n_11087);
  nand g27279 (n_9619, n_9955, n_11117);
  nand g27280 (n_9611, n_9910, n_11063);
  nand g27281 (n_9610, n_9914, n_11090);
  nand g27282 (n_9647, n_9886, n_11075);
  nand g27283 (n_9617, n_9915, n_11111);
  nand g27284 (n_9603, n_9889, n_11078);
  nand g27285 (n_12317, n_9573, n_9915);
  nand g27286 (n_9645, n_9585, n_11051);
  nand g27287 (n_9632, n_9924, n_11108);
  nand g27288 (n_9631, n_9961, n_11069);
  nand g27289 (n_11124, n_10005, n_10004);
  or g27290 (n_11117, wc232, n_9400);
  not gc232 (wc232, n_9551);
  or g27293 (n_12343, n_9317, wc233);
  not gc233 (wc233, n_9533);
  or g27298 (n_11102, wc234, b3);
  not gc234 (wc234, n_9548);
  or g27300 (n_11078, wc235, b8);
  not gc235 (wc235, n_9533);
  or g27301 (n_11072, wc236, b10);
  not gc236 (wc236, n_9527);
  or g27302 (n_11114, wc237, b1);
  not gc237 (wc237, n_9551);
  or g27303 (n_9528, n_9527, wc238);
  not gc238 (wc238, b9);
  or g27304 (n_11075, wc239, b9);
  not gc239 (wc239, n_9538);
  or g27305 (n_11084, wc240, b6);
  not gc240 (wc240, n_9567);
  or g27306 (n_11090, wc241, b5);
  not gc241 (wc241, n_9544);
  or g27307 (n_11105, wc242, b2);
  not gc242 (wc242, n_9555);
  or g27308 (n_11096, wc243, b4);
  not gc243 (wc243, n_9561);
  or g27309 (n_12756, wc244, b8);
  not gc244 (wc244, n_9538);
  or g27310 (n_12757, n_9538, wc245);
  not gc245 (wc245, b8);
  nand g27311 (n_9644, n_12756, n_12757);
  or g27312 (n_11111, wc246, b2);
  not gc246 (wc246, n_9551);
  or g27313 (n_11108, wc247, b3);
  not gc247 (wc247, n_9555);
  or g27314 (n_11099, wc248, b4);
  not gc248 (wc248, n_9548);
  or g27315 (n_11093, wc249, b5);
  not gc249 (wc249, n_9561);
  or g27316 (n_11087, wc250, b6);
  not gc250 (wc250, n_9544);
  or g27317 (n_11081, wc251, b7);
  not gc251 (wc251, n_9567);
  or g27318 (n_9567, n_10993, n_10994);
  or g27319 (n_9555, n_10957, n_10958);
  or g27320 (n_9533, n_11029, n_11030);
  or g27321 (n_9544, n_10975, n_10976);
  or g27322 (n_9548, n_11011, n_11012);
  nand g27323 (n_12758, n_9550, a6);
  or g27324 (n_12759, n_9550, a6);
  nand g27325 (n_9551, n_12758, n_12759);
  or g27327 (n_9561, n_11047, n_11048);
  or g27328 (n_9538, n_10939, n_10940);
  nand g27329 (n_11047, n_11043, n_11044);
  nand g27330 (n_11011, n_11007, n_11008);
  nand g27331 (n_11029, n_11025, n_11026);
  nand g27332 (n_10939, n_10935, n_10936);
  nand g27333 (n_10975, n_10971, n_10972);
  nand g27336 (n_10922, n_10919, n_10920);
  nand g27337 (n_10957, n_10953, n_10954);
  nand g27338 (n_10993, n_10989, n_10990);
  nand g27339 (n_11030, n_11027, n_11028);
  nand g27340 (n_10976, n_10973, n_10974);
  or g27341 (n_10004, n_9513, n_9378);
  nand g27345 (n_11125, n_9513, n_9378);
  nand g27347 (n_10940, n_10937, n_10938);
  nand g27348 (n_11048, n_11045, n_11046);
  nand g27350 (n_9952, n_9514, n_9524);
  nand g27351 (n_10994, n_10991, n_10992);
  nand g27353 (n_11012, n_11009, n_11010);
  nand g27354 (n_10958, n_10955, n_10956);
  nand g27357 (n_11028, n_9476, n_9512);
  nand g27358 (n_11046, n_9487, n_9512);
  or g27359 (n_9513, n_9459, wc252);
  not gc252 (wc252, n_9512);
  nand g27360 (n_10992, n_9493, n_9512);
  nand g27361 (n_10974, n_9480, n_9512);
  or g27362 (n_9514, wc253, n_9512);
  not gc253 (wc253, n_9501);
  nand g27363 (n_10938, n_9499, n_9512);
  nand g27364 (n_10956, n_9512, a7);
  nand g27365 (n_10921, n_9472, n_9512);
  nand g27366 (n_11010, n_9483, n_9512);
  or g27367 (n_11009, wc254, n_9525);
  not gc254 (wc254, n_10177);
  or g27368 (n_10991, wc255, n_9525);
  not gc255 (wc255, n_10168);
  or g27369 (n_11027, wc256, n_9525);
  not gc256 (wc256, n_10183);
  or g27370 (n_10973, wc257, n_9525);
  not gc257 (wc257, n_10162);
  or g27371 (n_10920, wc258, n_9525);
  not gc258 (wc258, n_10118);
  or g27372 (n_11045, wc259, n_9525);
  not gc259 (wc259, n_10201);
  or g27374 (n_10937, wc260, n_9525);
  not gc260 (wc260, n_10132);
  or g27375 (n_10955, wc261, n_9525);
  not gc261 (wc261, n_10153);
  nand g27384 (n_12260, n_12257, n_12258);
  or g27385 (n_9501, n_10907, b15);
  nand g27389 (n_9524, n_9369, n_10910);
  or g27390 (n_10907, n_10906, n_9321);
  or g27391 (n_12258, wc262, n_9459);
  not gc262 (wc262, n_10145);
  or g27393 (n_10910, wc263, n_9523);
  not gc263 (wc263, n_10125);
  or g27394 (n_10145, n_10886, wc264);
  not gc264 (wc264, b9);
  nand g27395 (n_10905, n_10902, n_10903);
  nand g27396 (n_10886, n_10885, n_9850);
  or g27397 (n_12257, n_10885, b9);
  or g27398 (n_10125, n_12197, n_9516);
  nand g27399 (n_12762, n_9515, n_9500);
  or g27400 (n_12763, n_9515, n_9500);
  nand g27401 (n_10118, n_12762, n_12763);
  nand g27402 (n_10885, n_9503, n_9511);
  nand g27403 (n_12764, n_9526, n_9511);
  or g27404 (n_12765, n_9526, n_9511);
  nand g27405 (n_10119, n_12764, n_12765);
  or g27406 (n_12197, n_12196, wc265);
  not gc265 (wc265, n_10829);
  nand g27408 (n_12196, n_12194, n_12195);
  nand g27409 (n_9500, n_10853, n_12221);
  nand g27410 (n_9511, n_10850, n_12218);
  nand g27411 (n_12218, n_9929, n_9510);
  nand g27413 (n_12766, n_9535, n_9522);
  or g27414 (n_12767, n_9535, n_9522);
  nand g27415 (n_10133, n_12766, n_12767);
  nand g27416 (n_12768, n_9536, n_9510);
  or g27417 (n_12769, n_9536, n_9510);
  nand g27418 (n_10134, n_12768, n_12769);
  nand g27419 (n_12770, n_9537, n_9495);
  or g27420 (n_12771, n_9537, n_9495);
  nand g27421 (n_10132, n_12770, n_12771);
  nand g27422 (n_12221, n_9930, n_9495);
  nand g27423 (n_9510, n_10844, n_12212);
  nand g27424 (n_9495, n_10847, n_12215);
  nand g27425 (n_9522, n_10835, n_12203);
  nand g27426 (n_12772, n_9530, n_9521);
  or g27427 (n_12773, n_9530, n_9521);
  nand g27428 (n_10184, n_12772, n_12773);
  nand g27429 (n_12215, n_9933, n_9494);
  nand g27430 (n_12203, n_9931, n_9521);
  nand g27431 (n_12774, n_9531, n_9509);
  or g27432 (n_12775, n_9531, n_9509);
  nand g27433 (n_10185, n_12774, n_12775);
  nand g27434 (n_12212, n_9906, n_9509);
  nand g27435 (n_12776, n_9532, n_9494);
  or g27436 (n_12777, n_9532, n_9494);
  nand g27437 (n_10183, n_12776, n_12777);
  nand g27438 (n_9509, n_10856, n_12224);
  nand g27439 (n_9521, n_10832, n_12200);
  nand g27440 (n_9494, n_10859, n_12227);
  nand g27441 (n_12778, n_9565, n_9508);
  or g27442 (n_12779, n_9565, n_9508);
  nand g27443 (n_10170, n_12778, n_12779);
  nand g27444 (n_12227, n_9935, n_9489);
  nand g27445 (n_12224, n_9934, n_9508);
  nand g27446 (n_12780, n_9566, n_9489);
  or g27447 (n_12781, n_9566, n_9489);
  nand g27448 (n_10168, n_12780, n_12781);
  nand g27449 (n_12200, n_9936, n_9520);
  nand g27450 (n_12782, n_9564, n_9520);
  or g27451 (n_12783, n_9564, n_9520);
  nand g27452 (n_10169, n_12782, n_12783);
  nand g27453 (n_9489, n_10862, n_12230);
  nand g27454 (n_9508, n_10865, n_12233);
  nand g27455 (n_9520, n_10838, n_12206);
  nand g27456 (n_12784, n_9543, n_9507);
  or g27457 (n_12785, n_9543, n_9507);
  nand g27458 (n_10164, n_12784, n_12785);
  nand g27459 (n_12206, n_9965, n_9519);
  nand g27460 (n_12233, n_9938, n_9507);
  nand g27461 (n_12786, n_9542, n_9519);
  or g27462 (n_12787, n_9542, n_9519);
  nand g27463 (n_10163, n_12786, n_12787);
  nand g27464 (n_12230, n_9939, n_9488);
  nand g27465 (n_12788, n_9541, n_9488);
  or g27466 (n_12789, n_9541, n_9488);
  nand g27467 (n_10162, n_12788, n_12789);
  nand g27468 (n_9507, n_10868, n_12236);
  nand g27469 (n_9488, n_10871, n_12239);
  nand g27470 (n_9519, n_10841, n_12209);
  nand g27471 (n_12236, n_9998, n_9506);
  nand g27472 (n_12239, n_9903, n_9484);
  nand g27473 (n_12790, n_9484, n_9560);
  or g27474 (n_12791, n_9484, n_9560);
  nand g27475 (n_10201, n_12790, n_12791);
  nand g27476 (n_12792, n_9559, n_9518);
  or g27477 (n_12793, n_9559, n_9518);
  nand g27478 (n_10202, n_12792, n_12793);
  nand g27479 (n_12794, n_9506, n_9558);
  or g27480 (n_12795, n_9506, n_9558);
  nand g27481 (n_10203, n_12794, n_12795);
  nand g27482 (n_12209, n_10002, n_9518);
  nand g27483 (n_9518, n_10874, n_12242);
  nand g27484 (n_12796, n_9505, n_9547);
  or g27485 (n_12797, n_9505, n_9547);
  nand g27486 (n_10179, n_12796, n_12797);
  nand g27487 (n_9484, n_10877, n_12245);
  or g27488 (n_12798, n_9481, n_9546);
  nand g27489 (n_12799, n_9481, n_9546);
  nand g27490 (n_10177, n_12798, n_12799);
  or g27491 (n_10904, n_10901, wc266);
  not gc266 (wc266, n_9459);
  nand g27492 (n_9506, n_10880, n_12248);
  nand g27493 (n_12800, n_9517, n_9545);
  or g27494 (n_12801, n_9517, n_9545);
  nand g27495 (n_10178, n_12800, n_12801);
  nand g27496 (n_9532, n_9933, n_10847);
  nand g27497 (n_9565, n_9934, n_10856);
  nand g27498 (n_10072, n_10825, n_10826);
  nand g27499 (n_9564, n_9936, n_10832);
  nand g27500 (n_9566, n_9935, n_10859);
  nand g27501 (n_9531, n_9906, n_10844);
  nand g27502 (n_9543, n_9938, n_10865);
  nand g27503 (n_9542, n_9965, n_10838);
  nand g27504 (n_9541, n_9939, n_10862);
  nand g27505 (n_9558, n_9998, n_10868);
  nand g27506 (n_9559, n_10002, n_10841);
  nand g27507 (n_9560, n_9903, n_10871);
  nand g27508 (n_9547, n_9967, n_10880);
  nand g27509 (n_9545, n_9986, n_10874);
  nand g27510 (n_9523, n_10819, n_10820);
  nand g27511 (n_12242, n_9517, n_9986);
  nand g27512 (n_12248, n_9505, n_9967);
  nand g27513 (n_10901, n_9850, n_9317);
  nand g27514 (n_9546, n_9984, n_10877);
  nand g27515 (n_12245, n_9481, n_9984);
  nand g27516 (n_9536, n_9929, n_10850);
  nand g27517 (n_9535, n_9869, n_10829);
  nand g27518 (n_9537, n_9930, n_10853);
  nand g27519 (n_9530, n_9931, n_10835);
  or g27520 (n_10880, wc267, b2);
  not gc267 (wc267, n_9483);
  or g27521 (n_10877, wc268, b1);
  not gc268 (wc268, n_9483);
  or g27522 (n_10903, n_9802, n_9472);
  or g27523 (n_10853, wc269, b6);
  not gc269 (wc269, n_9499);
  or g27524 (n_10862, wc270, b3);
  not gc270 (wc270, n_9480);
  or g27525 (n_10819, n_10817, wc271);
  not gc271 (wc271, n_9472);
  or g27526 (n_10856, wc272, b5);
  not gc272 (wc272, n_9493);
  or g27528 (n_12195, wc273, n_9472);
  not gc273 (wc273, n_9381);
  or g27529 (n_10871, wc274, b2);
  not gc274 (wc274, n_9487);
  or g27530 (n_12259, n_9328, wc275);
  not gc275 (wc275, n_9472);
  or g27531 (n_10874, wc276, n_9400);
  not gc276 (wc276, n_9483);
  or g27536 (n_10868, wc277, b3);
  not gc277 (wc277, n_9487);
  or g27537 (n_10859, wc278, b4);
  not gc278 (wc278, n_9493);
  or g27538 (n_12802, wc279, b7);
  not gc279 (wc279, n_9472);
  or g27539 (n_12803, n_9472, wc280);
  not gc280 (wc280, b7);
  nand g27540 (n_9515, n_12802, n_12803);
  or g27541 (n_10850, wc281, b7);
  not gc281 (wc281, n_9499);
  or g27542 (n_10847, wc282, b5);
  not gc282 (wc282, n_9476);
  or g27543 (n_10826, wc283, n_9472);
  not gc283 (wc283, n_9963);
  or g27544 (n_10844, wc284, b6);
  not gc284 (wc284, n_9476);
  or g27545 (n_10865, wc285, b4);
  not gc285 (wc285, n_9480);
  or g27546 (n_9480, n_10753, n_10754);
  nand g27547 (n_12804, n_9482, a8);
  or g27548 (n_12805, n_9482, a8);
  nand g27549 (n_9483, n_12804, n_12805);
  or g27551 (n_10817, n_9516, n_9381);
  or g27552 (n_9493, n_10807, n_10808);
  or g27553 (n_9499, n_10789, n_10790);
  or g27554 (n_9487, n_10735, n_10736);
  or g27555 (n_9476, n_10771, n_10772);
  nand g27556 (n_10808, n_10805, n_10806);
  or g27557 (n_10820, n_10818, n_9382);
  nand g27559 (n_10753, n_10749, n_10750);
  nand g27560 (n_10736, n_10733, n_10734);
  nand g27561 (n_10718, n_10715, n_10716);
  nand g27562 (n_10735, n_10731, n_10732);
  nand g27563 (n_10825, n_9317, n_9981);
  nand g27564 (n_10789, n_10785, n_10786);
  nand g27565 (n_10790, n_10787, n_10788);
  nand g27566 (n_10771, n_10767, n_10768);
  nand g27569 (n_10772, n_10769, n_10770);
  nand g27570 (n_10807, n_10803, n_10804);
  nand g27571 (n_10754, n_10751, n_10752);
  or g27572 (n_10805, wc286, n_9461);
  not gc286 (wc286, n_10192);
  or g27573 (n_10804, wc287, n_9471);
  not gc287 (wc287, n_10193);
  or g27574 (n_10769, wc288, n_9461);
  not gc288 (wc288, n_10186);
  or g27575 (n_10768, wc289, n_9471);
  not gc289 (wc289, n_10187);
  or g27576 (n_10787, wc290, n_9461);
  not gc290 (wc290, n_10189);
  or g27577 (n_10786, wc291, n_9471);
  not gc291 (wc291, n_10190);
  or g27578 (n_9963, n_9459, b8);
  or g27580 (n_10716, wc292, n_9461);
  not gc292 (wc292, n_10120);
  or g27581 (n_10733, wc293, n_9461);
  not gc293 (wc293, n_10147);
  or g27582 (n_10750, wc294, n_9471);
  not gc294 (wc294, n_10181);
  or g27584 (n_10751, wc295, n_9461);
  not gc295 (wc295, n_10180);
  nand g27585 (n_10706, n_9459, n_9382);
  or g27586 (n_10818, n_9379, n_9459);
  nand g27587 (n_9948, n_9470, n_9461);
  or g27588 (n_10732, wc296, n_9471);
  not gc296 (wc296, n_10148);
  nand g27589 (n_10752, n_9437, n_9458);
  nand g27590 (n_10806, n_9458, n_9441);
  nand g27591 (n_10788, n_9458, n_9447);
  nand g27593 (n_10734, n_9458, a9);
  nand g27596 (n_10717, n_9458, n_9428);
  nand g27599 (n_10770, n_9458, n_9434);
  or g27600 (n_9449, n_10694, n_9322);
  or g27601 (n_9458, n_10703, n_9333);
  nand g27602 (n_10694, n_10692, n_10693);
  nand g27603 (n_10703, n_10701, n_10702);
  or g27604 (n_10803, wc297, n_9470);
  not gc297 (wc297, n_10194);
  or g27605 (n_10749, wc298, n_9470);
  not gc298 (wc298, n_10182);
  nand g27606 (n_10702, n_10116, n_9419);
  nand g27607 (n_10693, n_10066, n_9419);
  or g27608 (n_10767, wc299, n_9470);
  not gc299 (wc299, n_10188);
  or g27609 (n_10731, wc300, n_9470);
  not gc300 (wc300, n_10149);
  or g27610 (n_10785, wc301, n_9470);
  not gc301 (wc301, n_10191);
  nand g27611 (n_10692, n_10673, b6);
  or g27612 (n_10066, n_10673, b6);
  nand g27614 (n_10701, n_10682, b7);
  or g27615 (n_10116, n_10682, b7);
  nand g27616 (n_10682, n_10680, n_10604);
  nand g27617 (n_10673, n_10672, n_9430);
  nand g27618 (n_10685, n_10094, n_9465);
  or g27619 (n_10680, wc302, n_9457);
  not gc302 (wc302, n_9451);
  or g27620 (n_10672, wc303, n_9448);
  not gc303 (wc303, n_9429);
  nand g27621 (n_12808, n_9460, n_9457);
  or g27622 (n_12809, n_9460, n_9457);
  nand g27623 (n_10120, n_12808, n_12809);
  nand g27624 (n_9465, n_10654, n_10655);
  nand g27628 (n_10655, n_10018, n_9419);
  nand g27629 (n_9457, n_10616, n_12164);
  nand g27630 (n_9448, n_10613, n_12161);
  or g27631 (n_10018, n_10649, n_9355);
  nand g27632 (n_10654, n_10649, n_9355);
  or g27633 (n_10094, n_10667, wc304);
  not gc304 (wc304, n_9462);
  nand g27634 (n_12164, n_9909, n_9456);
  nand g27635 (n_12161, n_9970, n_9443);
  nand g27636 (n_12812, n_9861, n_9496);
  or g27637 (n_12813, n_9861, n_9496);
  nand g27638 (n_10191, n_12812, n_12813);
  nand g27639 (n_12814, n_9497, n_9443);
  or g27640 (n_12815, n_9497, n_9443);
  nand g27641 (n_10190, n_12814, n_12815);
  nand g27642 (n_12816, n_9498, n_9456);
  or g27643 (n_12817, n_9498, n_9456);
  nand g27644 (n_10189, n_12816, n_12817);
  nand g27645 (n_9443, n_10622, n_12170);
  nand g27646 (n_9456, n_10619, n_12167);
  nand g27647 (n_10649, n_10647, n_10648);
  or g27648 (n_10667, n_10666, n_9469);
  nand g27649 (n_12818, n_9475, n_9468);
  or g27650 (n_12819, n_9475, n_9468);
  nand g27651 (n_10188, n_12818, n_12819);
  nand g27652 (n_12167, n_9896, n_9455);
  nand g27653 (n_10647, n_9352, n_9887);
  nand g27654 (n_9469, n_10607, n_9468);
  nand g27655 (n_12820, n_9474, n_9442);
  or g27656 (n_12821, n_9474, n_9442);
  nand g27657 (n_10187, n_12820, n_12821);
  nand g27658 (n_12170, n_9898, n_9442);
  nand g27659 (n_12822, n_9473, n_9455);
  or g27660 (n_12823, n_9473, n_9455);
  nand g27661 (n_10186, n_12822, n_12823);
  or g27662 (n_10648, wc305, n_9428);
  not gc305 (wc305, n_9464);
  nand g27663 (n_9442, n_10628, n_12176);
  nand g27664 (n_9468, n_10610, n_12158);
  nand g27665 (n_9455, n_10625, n_12173);
  nand g27666 (n_12158, n_9900, n_9467);
  nand g27667 (n_9464, n_9462, n_10631);
  nand g27668 (n_12824, n_9454, n_9490);
  or g27669 (n_12825, n_9454, n_9490);
  nand g27670 (n_10192, n_12824, n_12825);
  nand g27671 (n_12173, n_9917, n_9454);
  nand g27672 (n_12826, n_9492, n_9467);
  or g27673 (n_12827, n_9492, n_9467);
  nand g27674 (n_10194, n_12826, n_12827);
  nand g27675 (n_12828, n_9438, n_9491);
  or g27676 (n_12829, n_9438, n_9491);
  nand g27677 (n_10193, n_12828, n_12829);
  nand g27678 (n_12176, n_9951, n_9438);
  nand g27679 (n_9467, n_10634, n_12179);
  nand g27680 (n_9475, n_9463, n_10607);
  nand g27681 (n_9490, n_9917, n_10625);
  nand g27682 (n_12830, n_9453, n_9479);
  or g27683 (n_12831, n_9453, n_9479);
  nand g27684 (n_10180, n_12830, n_12831);
  nand g27685 (n_9496, n_9462, n_9944);
  nand g27686 (n_9491, n_9951, n_10628);
  or g27687 (n_12832, n_9435, n_9478);
  nand g27688 (n_12833, n_9435, n_9478);
  nand g27689 (n_10181, n_12832, n_12833);
  nand g27690 (n_9492, n_9900, n_10610);
  nand g27691 (n_9438, n_10637, n_12182);
  nand g27692 (n_9460, n_9451, n_10604);
  nand g27693 (n_9498, n_9909, n_10616);
  nand g27694 (n_10631, n_9463, n_9944);
  nand g27695 (n_9454, n_10640, n_12185);
  nand g27696 (n_9473, n_9896, n_10619);
  nand g27697 (n_9474, n_9898, n_10622);
  nand g27698 (n_12834, n_9466, n_9477);
  or g27699 (n_12835, n_9466, n_9477);
  nand g27700 (n_10182, n_12834, n_12835);
  nand g27701 (n_10666, n_10664, n_10665);
  nand g27702 (n_9497, n_9970, n_10613);
  or g27703 (n_10619, wc306, b4);
  not gc306 (wc306, n_9434);
  or g27704 (n_10622, wc307, b3);
  not gc307 (wc307, n_9434);
  nand g27705 (n_12179, n_9466, n_10003);
  nand g27707 (n_12185, n_9453, n_9919);
  nand g27709 (n_9477, n_10003, n_10634);
  or g27710 (n_10665, wc308, n_9428);
  not gc308 (wc308, n_9352);
  or g27712 (n_10628, wc309, b2);
  not gc309 (wc309, n_9441);
  or g27713 (n_10613, wc310, b4);
  not gc310 (wc310, n_9447);
  nand g27714 (n_9478, n_9920, n_10637);
  nand g27715 (n_9479, n_9919, n_10640);
  nand g27716 (n_12182, n_9435, n_9920);
  or g27717 (n_10604, n_9428, wc311);
  not gc311 (wc311, b6);
  or g27718 (n_10625, wc312, b3);
  not gc312 (wc312, n_9441);
  or g27719 (n_10616, wc313, b5);
  not gc313 (wc313, n_9447);
  or g27721 (n_9434, n_10588, n_10589);
  or g27722 (n_9441, n_10570, n_10571);
  or g27723 (n_9447, n_10552, n_10553);
  or g27724 (n_10640, wc314, b2);
  not gc314 (wc314, n_9437);
  or g27725 (n_10634, wc315, n_9400);
  not gc315 (wc315, n_9437);
  or g27726 (n_10637, wc316, b1);
  not gc316 (wc316, n_9437);
  nand g27727 (n_10588, n_10584, n_10585);
  nand g27728 (n_10570, n_10566, n_10567);
  nand g27729 (n_12836, n_9436, a10);
  or g27730 (n_12837, n_9436, a10);
  nand g27731 (n_9437, n_12836, n_12837);
  nand g27732 (n_10552, n_10548, n_10549);
  nand g27733 (n_10601, n_10598, n_10599);
  or g27734 (n_10584, wc317, n_9426);
  not gc317 (wc317, n_10197);
  or g27738 (n_10566, wc318, n_9426);
  not gc318 (wc318, n_10158);
  or g27739 (n_10548, wc319, n_9426);
  not gc319 (wc319, n_10140);
  nand g27740 (n_10553, n_10550, n_10551);
  nand g27742 (n_10589, n_10586, n_10587);
  nand g27744 (n_9918, n_9425, n_9420);
  nand g27745 (n_10571, n_10568, n_10569);
  or g27748 (n_9425, n_10535, n_9352);
  nand g27752 (n_10664, n_9419, n_9355);
  nand g27754 (n_10569, n_9418, a11);
  nand g27755 (n_10587, n_9406, n_9418);
  nand g27757 (n_10600, n_9402, n_9418);
  or g27758 (n_9420, n_9418, wc320);
  not gc320 (wc320, n_9411);
  or g27759 (n_10535, n_10534, n_9355);
  nand g27760 (n_10551, n_9409, n_9418);
  or g27763 (n_9418, n_12131, n_10283);
  or g27764 (n_10534, n_10533, n_9383);
  or g27765 (n_9411, n_10517, n_9323);
  or g27766 (n_10517, n_10515, n_10516);
  nand g27767 (n_10533, n_10531, n_10532);
  or g27768 (n_12131, n_12129, n_12130);
  nand g27769 (n_10516, n_10513, n_10514);
  or g27770 (n_10532, wc321, n_10530);
  not gc321 (wc321, n_9424);
  nand g27771 (n_12130, n_12127, n_12128);
  or g27775 (n_10514, n_10510, n_9410);
  nand g27776 (n_12842, n_9421, n_9417);
  or g27777 (n_12843, n_9421, n_9417);
  nand g27778 (n_10123, n_12842, n_12843);
  or g27779 (n_12128, n_12124, n_9417);
  or g27780 (n_9424, n_12140, wc322);
  not gc322 (wc322, n_10478);
  nand g27781 (n_12140, n_12138, n_12139);
  nand g27782 (n_9417, n_10484, n_12146);
  nand g27783 (n_9410, n_10481, n_12143);
  nand g27784 (n_12146, n_9972, n_9416);
  nand g27786 (n_12844, n_9444, n_9407);
  or g27787 (n_12845, n_9444, n_9407);
  nand g27788 (n_10140, n_12844, n_12845);
  nand g27789 (n_12846, n_9445, n_9416);
  or g27790 (n_12847, n_9445, n_9416);
  nand g27791 (n_10138, n_12846, n_12847);
  nand g27792 (n_12143, n_9973, n_9407);
  nand g27793 (n_12848, n_9446, n_9423);
  or g27794 (n_12849, n_9446, n_9423);
  nand g27795 (n_10139, n_12848, n_12849);
  nand g27796 (n_9444, n_9973, n_10481);
  or g27797 (n_12850, n_9404, n_9432);
  nand g27798 (n_12851, n_9404, n_9432);
  nand g27799 (n_10197, n_12850, n_12851);
  nand g27800 (n_12852, n_9422, n_9431);
  or g27801 (n_12853, n_9422, n_9431);
  nand g27802 (n_10196, n_12852, n_12853);
  nand g27803 (n_12854, n_9415, n_9433);
  or g27804 (n_12855, n_9415, n_9433);
  nand g27805 (n_10195, n_12854, n_12855);
  nand g27806 (n_9445, n_9972, n_10484);
  nand g27807 (n_9446, n_9932, n_10478);
  nand g27808 (n_9423, n_10487, n_12149);
  nand g27809 (n_9407, n_10490, n_12152);
  nand g27810 (n_9416, n_10493, n_12155);
  nand g27812 (n_12152, n_9404, n_9977);
  nand g27813 (n_12129, n_12125, n_12126);
  or g27814 (n_12127, n_9817, wc323);
  not gc323 (wc323, b4);
  nand g27815 (n_9432, n_9977, n_10490);
  nand g27817 (n_10515, n_10511, n_10512);
  nand g27818 (n_9431, n_9975, n_10487);
  or g27819 (n_10513, n_9817, wc324);
  not gc324 (wc324, b3);
  nand g27820 (n_12124, n_9921, n_9413);
  or g27821 (n_10481, wc325, b2);
  not gc325 (wc325, n_9409);
  or g27822 (n_10484, wc326, b3);
  not gc326 (wc326, n_9409);
  nand g27823 (n_9433, n_9912, n_10493);
  nand g27824 (n_10510, n_10070, n_9403);
  nand g27825 (n_9421, n_9413, n_10472);
  nand g27826 (n_12149, n_9422, n_9975);
  nand g27827 (n_12155, n_9415, n_9912);
  nand g27828 (n_10530, n_10079, n_10078);
  or g27829 (n_12138, wc327, n_9402);
  not gc327 (wc327, n_9346);
  or g27830 (n_9409, n_10468, n_10469);
  or g27832 (n_10511, n_9800, n_9402);
  or g27833 (n_10490, wc328, b1);
  not gc328 (wc328, n_9406);
  or g27834 (n_12125, n_9347, n_9402);
  or g27835 (n_9817, wc329, n_9402);
  not gc329 (wc329, n_9393);
  or g27836 (n_10493, wc330, b2);
  not gc330 (wc330, n_9406);
  or g27837 (n_10487, wc331, n_9400);
  not gc331 (wc331, n_9406);
  or g27838 (n_10472, n_9402, wc332);
  not gc332 (wc332, b4);
  nand g27839 (n_10468, n_9809, n_10465);
  nand g27840 (n_12856, n_9405, a12);
  or g27841 (n_12857, n_9405, a12);
  nand g27842 (n_9406, n_12856, n_12857);
  nand g27846 (n_10465, n_10161, a13);
  nand g27847 (n_10469, n_10466, n_10467);
  nand g27848 (n_10454, n_10451, n_10452);
  or g27849 (n_10070, n_9393, b4);
  or g27850 (n_10451, wc333, n_9394);
  not gc333 (wc333, n_10144);
  nand g27851 (n_12126, n_9393, b5);
  or g27852 (n_9921, n_9393, b5);
  or g27853 (n_10467, wc334, n_9394);
  not gc334 (wc334, n_10159);
  nand g27854 (n_10531, n_9393, n_9349);
  nand g27855 (n_10512, n_9393, b4);
  or g27856 (n_10078, n_9393, n_9349);
  nand g27858 (n_9941, n_9394, n_9401);
  or g27860 (n_10439, n_9816, b0);
  or g27861 (n_9809, n_9816, n_9337);
  or g27864 (n_10453, n_10450, n_9816);
  or g27868 (n_9392, n_10436, n_9334);
  or g27869 (n_9387, n_10427, n_9315);
  nand g27870 (n_10436, n_10434, n_10435);
  or g27872 (n_10427, n_10426, n_9323);
  or g27873 (n_9401, n_10394, n_9383);
  nand g27874 (n_10435, n_10074, n_9341);
  or g27875 (n_10394, n_10393, n_9356);
  or g27876 (n_10426, wc335, n_10425);
  not gc335 (wc335, n_10424);
  or g27877 (n_10074, n_10406, b3);
  nand g27878 (n_10434, n_10406, b3);
  or g27879 (n_10424, n_10421, n_9337);
  or g27880 (n_10393, n_10391, n_10392);
  nand g27881 (n_10406, n_10404, n_10397);
  nand g27882 (n_12860, n_9396, n_9391);
  or g27883 (n_12861, n_9396, n_9391);
  nand g27884 (n_10144, n_12860, n_12861);
  nand g27885 (n_10391, n_10387, n_10388);
  nand g27886 (n_10425, n_10422, n_10423);
  or g27887 (n_10404, wc336, n_9391);
  not gc336 (wc336, n_9389);
  nand g27888 (n_9396, n_9389, n_10397);
  nand g27889 (n_10421, n_9947, n_9386);
  or g27890 (n_10450, n_9386, wc337);
  not gc337 (wc337, n_9337);
  or g27891 (n_9389, n_9385, b2);
  nand g27892 (n_10397, n_9385, b2);
  nand g27893 (n_10388, n_9385, n_9400);
  or g27894 (n_9386, n_9385, b1);
  nand g27895 (n_10422, n_10073, n_9385);
  nand g27896 (n_9385, n_10092, a14);
  nand g27899 (n_9384, n_10369, n_10370);
  or g27900 (n_10370, n_10368, n_9357);
  or g27901 (n_10368, n_10367, n_9383);
  or g27902 (n_9383, n_10358, n_9382);
  or g27903 (n_10358, n_10357, n_9381);
  or g27904 (n_10357, n_9379, wc338);
  not gc338 (wc338, n_9369);
  or g27905 (n_9379, n_10352, n_9378);
  or g27906 (n_10352, n_9375, n_9377);
  or g27907 (n_9375, n_10349, n_9373);
  nand g27908 (n_9369, n_9331, n_9368);
  or g27909 (n_10349, n_10348, n_9372);
  or g27910 (n_12863, wc339, n_9331);
  not gc339 (wc339, n_9368);
  or g27911 (n_12864, n_9368, wc340);
  not gc340 (wc340, n_9331);
  nand g27912 (n_9373, n_12863, n_12864);
  or g27913 (n_9368, n_10343, wc341);
  not gc341 (wc341, n_9358);
  or g27914 (n_10348, n_9374, n_9371);
  or g27915 (n_12865, wc342, n_9318);
  not gc342 (wc342, n_9945);
  or g27916 (n_12866, n_9945, wc343);
  not gc343 (wc343, n_9318);
  nand g27917 (n_9374, n_12865, n_12866);
  nand g27918 (n_10343, n_10341, n_10342);
  nand g27919 (n_9945, n_9358, n_9367);
  or g27920 (n_10341, wc344, n_9367);
  not gc344 (wc344, n_9318);
  nand g27924 (n_9372, n_12867, n_12868);
  nand g27925 (n_9366, n_10057, n_9329);
  nand g27926 (n_9378, n_10333, n_10334);
  nand g27927 (n_10057, n_9360, n_10328);
  nand g27928 (n_12869, n_9894, n_9370);
  or g27929 (n_12870, n_9894, n_9370);
  nand g27930 (n_9371, n_12869, n_12870);
  nand g27932 (n_10328, n_9319, n_9880);
  nand g27933 (n_9370, n_9359, n_10325);
  nand g27934 (n_10325, n_9329, n_9365);
  nand g27935 (n_10333, n_10093, n_9365);
  or g27936 (n_9365, n_10322, wc345);
  not gc345 (wc345, n_9361);
  nand g27937 (n_10322, n_10321, n_9807);
  nand g27938 (n_12871, n_9968, n_9376);
  or g27939 (n_12872, n_9968, n_9376);
  nand g27940 (n_9377, n_12871, n_12872);
  or g27941 (n_10321, wc346, n_9364);
  not gc346 (wc346, n_9320);
  nand g27942 (n_9968, n_9361, n_9364);
  nand g27943 (n_9364, n_9328, n_9363);
  or g27944 (n_10367, n_9356, n_9925);
  nand g27945 (n_12873, n_9956, n_9363);
  or g27946 (n_12874, n_9956, n_9363);
  nand g27947 (n_9382, n_12873, n_12874);
  or g27948 (n_9356, n_10289, n_9352);
  or g27949 (n_9363, n_10295, wc347);
  not gc347 (wc347, n_9802);
  nand g27950 (n_12875, n_9905, n_9380);
  or g27951 (n_12876, n_9905, n_9380);
  nand g27952 (n_9381, n_12875, n_12876);
  nand g27953 (n_10295, n_10294, n_9353);
  or g27954 (n_10289, n_10288, n_9349);
  or g27955 (n_10288, n_9346, n_9355);
  or g27956 (n_10294, wc348, n_9362);
  not gc348 (wc348, n_9317);
  nand g27957 (n_10073, n_9808, n_10316);
  nand g27958 (n_10392, n_10389, n_10390);
  nand g27959 (n_12877, n_9987, n_9354);
  or g27960 (n_12878, n_9987, n_9354);
  nand g27961 (n_9355, n_12877, n_12878);
  nand g27962 (n_9362, n_9327, n_9354);
  nand g27963 (n_10389, n_9341, n_9357);
  or g27964 (n_10369, wc349, n_9340);
  not gc349 (wc349, n_9325);
  nand g27965 (n_10423, n_9341, b2);
  nand g27966 (n_10316, n_9341, b1);
  or g27970 (n_9947, n_9341, b2);
  or g27971 (n_9335, n_10313, b3);
  or g27972 (n_9325, n_10280, wc350);
  not gc350 (wc350, a15);
  nand g27973 (n_12880, n_9350, n_9351);
  or g27974 (n_12881, n_9350, n_9351);
  nand g27975 (n_9352, n_12880, n_12881);
  nand g27976 (n_9341, n_9340, a15);
  nand g27977 (n_12107, n_12106, n_9801);
  or g27978 (n_9340, n_10307, n_9338);
  nand g27980 (n_9350, n_9347, n_10274);
  or g27981 (n_10313, n_10312, b0);
  or g27982 (n_10280, n_10279, n_9315);
  or g27983 (n_10279, n_9323, n_9324);
  or g27984 (n_10307, n_10306, n_9334);
  nand g27985 (n_12882, n_9971, n_9348);
  or g27986 (n_12883, n_9971, n_9348);
  nand g27987 (n_9349, n_12882, n_12883);
  nand g27988 (n_10274, n_9326, n_9348);
  or g27989 (n_10312, n_9324, n_9334);
  or g27990 (n_9348, n_12086, wc351);
  not gc351 (wc351, n_9800);
  or g27991 (n_9334, n_10283, n_9326);
  or g27992 (n_9322, n_10241, b15);
  nand g27993 (n_12086, n_12085, n_9343);
  nand g27994 (n_12884, n_9344, n_9345);
  or g27995 (n_12885, n_9344, n_9345);
  nand g27996 (n_9346, n_12884, n_12885);
  or g27997 (n_10283, n_9333, n_9327);
  or g27998 (n_10241, n_9321, n_9317);
  or g27999 (n_12085, n_10238, wc352);
  not gc352 (wc352, n_9315);
  nand g28000 (n_9415, n_10246, n_10247);
  nand g28001 (n_9670, n_10270, n_10271);
  nand g28002 (n_9422, n_10247, n_12089);
  nand g28003 (n_9654, n_10271, n_12101);
  nand g28004 (n_9589, n_10265, n_12098);
  nand g28005 (n_9573, n_10264, n_10265);
  nand g28006 (n_10306, n_10304, n_10305);
  nand g28007 (n_9344, n_9343, n_10238);
  or g28008 (n_9333, n_9846, n_9328);
  nand g28009 (n_11860, n_11856, n_11857);
  nand g28010 (n_9466, n_10253, n_12092);
  nand g28011 (n_9517, n_10259, n_12095);
  nand g28012 (n_9505, n_10258, n_10259);
  nand g28013 (n_9453, n_10252, n_10253);
  nand g28014 (n_12886, n_9653, n_9747);
  or g28015 (n_12887, n_9653, n_9747);
  nand g28016 (n_10084, n_12886, n_12887);
  or g28017 (n_10252, wc353, b1);
  not gc353 (wc353, n_9864);
  nand g28018 (n_10238, n_9338, n_9342);
  or g28020 (n_10246, wc354, b1);
  not gc354 (wc354, n_9856);
  or g28021 (n_9846, n_9332, n_9329);
  nand g28022 (n_12888, n_9452, n_9486);
  or g28023 (n_12889, n_9452, n_9486);
  nand g28024 (n_10149, n_12888, n_12889);
  or g28025 (n_12101, wc355, b1);
  not gc355 (wc355, n_9862);
  or g28026 (n_10264, wc356, b1);
  not gc356 (wc356, n_9879);
  nand g28027 (n_12890, n_9974, n_9342);
  or g28028 (n_12891, n_9974, n_9342);
  nand g28029 (n_9357, n_12890, n_12891);
  nand g28030 (n_12433, n_9397, n_9768);
  nand g28032 (n_12892, n_9390, n_9408);
  or g28033 (n_12893, n_9390, n_9408);
  nand g28034 (n_10159, n_12892, n_12893);
  or g28036 (n_10258, wc357, b1);
  not gc357 (wc357, n_9875);
  or g28037 (n_12894, wc358, n_9399);
  not gc358 (wc358, n_9871);
  or g28038 (n_12895, n_9871, wc359);
  not gc359 (wc359, n_9399);
  nand g28039 (n_9400, n_12894, n_12895);
  nand g28041 (n_10304, n_9925, b1);
  or g28043 (n_12896, wc360, n_9398);
  not gc360 (wc360, n_9390);
  nand g28046 (n_9391, n_10217, n_12080);
  or g28047 (n_9321, n_10235, n_9319);
  nand g28048 (n_12898, n_9572, n_9626);
  or g28049 (n_12899, n_9572, n_9626);
  nand g28050 (n_10151, n_12898, n_12899);
  nand g28051 (n_12900, n_9504, n_9554);
  or g28052 (n_12901, n_9504, n_9554);
  nand g28053 (n_10154, n_12900, n_12901);
  nand g28054 (n_11856, n_9768, b1);
  nand g28055 (n_12902, n_9414, n_9440);
  or g28056 (n_12903, n_9414, n_9440);
  nand g28057 (n_10157, n_12902, n_12903);
  or g28058 (n_10387, n_9390, wc361);
  not gc361 (wc361, n_9398);
  nand g28059 (n_10253, n_9452, a9);
  or g28060 (n_12904, wc362, a9);
  not gc362 (wc362, n_9397);
  or g28061 (n_12905, n_9397, wc363);
  not gc363 (wc363, a9);
  nand g28062 (n_9486, n_12904, n_12905);
  nand g28063 (n_10148, n_9435, n_10223);
  nand g28064 (n_12906, n_9452, n_9485);
  or g28065 (n_12907, n_9452, n_9485);
  nand g28066 (n_10147, n_12906, n_12907);
  nand g28067 (n_9974, n_9338, n_9343);
  nand g28068 (n_9956, n_9328, n_9361);
  nand g28069 (n_10259, n_9504, a7);
  nand g28070 (n_9380, n_9317, n_9802);
  nand g28071 (n_12908, n_9414, n_9439);
  or g28072 (n_12909, n_9414, n_9439);
  nand g28073 (n_10156, n_12908, n_12909);
  or g28074 (n_10305, n_9339, a15);
  nand g28075 (n_12910, n_9504, n_9553);
  or g28076 (n_12911, n_9504, n_9553);
  nand g28077 (n_10155, n_12910, n_12911);
  or g28078 (n_12912, wc364, a7);
  not gc364 (wc364, n_9397);
  or g28079 (n_12913, n_9397, wc365);
  not gc365 (wc365, a7);
  nand g28080 (n_9554, n_12912, n_12913);
  or g28081 (n_10235, n_9320, n_9318);
  nand g28082 (n_10093, n_9359, n_9329);
  nand g28083 (n_10153, n_9481, n_10229);
  nand g28084 (n_9376, n_9320, n_9807);
  or g28085 (n_12914, wc366, a11);
  not gc366 (wc366, n_9397);
  or g28086 (n_12915, n_9397, wc367);
  not gc367 (wc367, a11);
  nand g28087 (n_9440, n_12914, n_12915);
  nand g28088 (n_10265, n_9572, a5);
  nand g28089 (n_10158, n_9404, n_10232);
  nand g28090 (n_9342, n_9808, n_9871);
  nand g28091 (n_9959, n_9330, n_9358);
  or g28092 (n_9332, n_9330, n_9331);
  nand g28093 (n_12916, n_9572, n_9625);
  or g28094 (n_12917, n_9572, n_9625);
  nand g28095 (n_10152, n_12916, n_12917);
  or g28096 (n_12918, wc368, a5);
  not gc368 (wc368, n_9397);
  or g28097 (n_12919, n_9397, wc369);
  not gc369 (wc369, a5);
  nand g28098 (n_9626, n_12918, n_12919);
  nand g28099 (n_10150, n_9549, n_10226);
  nand g28100 (n_10271, n_9653, a3);
  nand g28101 (n_9399, n_9324, n_9808);
  nand g28102 (n_9345, n_9800, n_9315);
  or g28103 (n_10390, wc370, a13);
  not gc370 (wc370, n_9397);
  nand g28104 (n_10247, n_9414, a11);
  nand g28105 (n_12920, n_9653, n_9746);
  or g28106 (n_12921, n_9653, n_9746);
  nand g28107 (n_10085, n_12920, n_12921);
  nand g28108 (n_9987, n_9327, n_9353);
  or g28109 (n_12922, wc371, a3);
  not gc371 (wc371, n_9397);
  or g28110 (n_12923, n_9397, wc372);
  not gc372 (wc372, a3);
  nand g28111 (n_9747, n_12922, n_12923);
  nand g28112 (n_9408, n_10000, n_10217);
  nand g28113 (n_10083, n_9621, n_10220);
  nand g28114 (n_9768, n_10214, a1);
  nand g28115 (n_9351, n_9316, n_9801);
  nand g28116 (n_9971, n_9347, n_9326);
  or g28117 (n_11857, n_9743, a0);
  nand g28118 (n_12080, n_9390, n_10000);
  nand g28119 (n_9801, b5, b6);
  nand g28120 (n_9358, b12, b13);
  nand g28121 (n_9802, b8, b7);
  nand g28122 (n_9807, b9, b10);
  nand g28123 (n_9800, b4, b3);
  nand g28124 (n_9361, b8, b9);
  nand g28125 (n_10342, b14, b13);
  or g28126 (n_9337, a13, wc373);
  not gc373 (wc373, b0);
  nand g28127 (n_9808, b2, b1);
  nand g28130 (n_9397, n_12924, n_12925);
  or g28131 (n_10217, wc374, b1);
  not gc374 (wc374, a13);
  or g28132 (n_9338, b2, b3);
  or g28133 (n_9404, a11, wc375);
  not gc375 (wc375, b0);
  or g28134 (n_10232, wc376, b0);
  not gc376 (wc376, a11);
  or g28135 (n_12926, wc377, b1);
  not gc377 (wc377, a11);
  or g28136 (n_12927, a11, wc378);
  not gc378 (wc378, b1);
  nand g28137 (n_9439, n_12926, n_12927);
  or g28138 (n_9435, a9, wc379);
  not gc379 (wc379, b0);
  or g28139 (n_10223, wc380, b0);
  not gc380 (wc380, a9);
  or g28140 (n_12928, wc381, b1);
  not gc381 (wc381, a9);
  or g28141 (n_12929, a9, wc382);
  not gc382 (wc382, b1);
  nand g28142 (n_9485, n_12928, n_12929);
  or g28143 (n_9481, a7, wc383);
  not gc383 (wc383, b0);
  or g28144 (n_9326, b4, b5);
  or g28145 (n_12930, wc384, b1);
  not gc384 (wc384, a7);
  or g28146 (n_12931, a7, wc385);
  not gc385 (wc385, b1);
  nand g28147 (n_9553, n_12930, n_12931);
  or g28148 (n_9327, b6, b7);
  or g28149 (n_10229, wc386, b0);
  not gc386 (wc386, a7);
  or g28150 (n_9328, b8, b9);
  or g28151 (n_9549, a5, wc387);
  not gc387 (wc387, b0);
  or g28152 (n_9329, b11, b10);
  or g28153 (n_9331, b14, b15);
  or g28154 (n_9330, b13, b12);
  or g28155 (n_12932, wc388, b1);
  not gc388 (wc388, a5);
  or g28156 (n_12933, a5, wc389);
  not gc389 (wc389, b1);
  nand g28157 (n_9625, n_12932, n_12933);
  or g28158 (n_10226, wc390, b0);
  not gc390 (wc390, a5);
  or g28159 (n_9315, b3, b4);
  or g28160 (n_9621, a3, wc391);
  not gc391 (wc391, b0);
  or g28161 (n_12934, wc392, b1);
  not gc392 (wc392, a3);
  or g28162 (n_12935, a3, wc393);
  not gc393 (wc393, b1);
  nand g28163 (n_9746, n_12934, n_12935);
  or g28164 (n_10220, wc394, b0);
  not gc394 (wc394, a3);
  or g28165 (n_10214, a0, wc395);
  not gc395 (wc395, b0);
  or g28166 (n_9318, b13, b14);
  and g28168 (o14, n_9335, n_9384);
  and g28169 (o13, n_9335, wc396);
  not gc396 (wc396, n_9387);
  and g28170 (o12, n_9335, n_9941);
  and g28171 (o11, n_9335, wc397);
  not gc397 (wc397, n_9411);
  and g28172 (o10, n_9335, n_9918);
  and g28173 (o9, n_9335, wc398);
  not gc398 (wc398, n_9449);
  and g28174 (o8, n_9335, n_9948);
  and g28175 (o7, n_9335, wc399);
  not gc399 (wc399, n_9501);
  and g28176 (o6, n_9335, n_9952);
  and g28177 (o5, n_9335, wc400);
  not gc400 (wc400, n_9570);
  and g28178 (o4, n_9335, n_9904);
  and g28179 (o3, n_9335, wc401);
  not gc401 (wc401, n_9650);
  and g28180 (o2, n_9335, n_9744);
  and g28182 (o0, n_10006, n_9335);
  or g28184 (n_12924, wc402, b1);
  not gc402 (wc402, b0);
  or g28185 (n_12925, b0, wc403);
  not gc403 (wc403, b1);
  or g28186 (n_12089, n_9397, wc404);
  not gc404 (wc404, n_9856);
  or g28187 (n_12092, n_9397, wc405);
  not gc405 (wc405, n_9864);
  or g28188 (n_12095, n_9397, wc406);
  not gc406 (wc406, n_9875);
  or g28189 (n_12098, n_9397, wc407);
  not gc407 (wc407, n_9879);
  or g28190 (n_10270, n_9397, wc408);
  not gc408 (wc408, n_9862);
  or g28192 (n_12106, n_10274, wc409);
  not gc409 (wc409, n_9316);
  or g28193 (n_9354, n_12107, wc410);
  not gc410 (wc410, n_9347);
  and g28194 (o15, wc411, n_9335);
  not gc411 (wc411, n_9325);
  or g28195 (n_10334, wc412, n_9880);
  not gc412 (wc412, n_9329);
  or g28196 (n_9367, wc413, n_9366);
  not gc413 (wc413, n_9330);
  or g28197 (n_12867, wc414, n_9366);
  not gc414 (wc414, n_9959);
  or g28198 (n_12868, n_9959, wc415);
  not gc415 (wc415, n_9366);
  or g28199 (n_10466, n_9401, n_12896);
  or g28200 (n_9816, wc416, n_9387);
  not gc416 (wc416, n_9401);
  or g28201 (n_9394, wc417, n_9392);
  not gc417 (wc417, n_9387);
  or g28202 (n_10452, n_9385, wc418);
  not gc418 (wc418, n_9392);
  or g28203 (n_9393, n_9341, wc419);
  not gc419 (wc419, n_9392);
  or g28204 (n_10161, n_9392, wc420);
  not gc420 (wc420, n_10439);
  or g28205 (n_9402, wc421, n_10454);
  not gc421 (wc421, n_10453);
  or g28207 (n_9932, n_9357, wc422);
  not gc422 (wc422, n_9409);
  or g28208 (n_10478, wc423, n_9409);
  not gc423 (wc423, n_9357);
  or g28209 (n_12139, wc424, n_9423);
  not gc424 (wc424, n_9932);
  or g28210 (n_12840, wc425, n_9403);
  not gc425 (wc425, n_9410);
  or g28212 (n_9419, n_9393, wc426);
  not gc426 (wc426, n_9418);
  or g28213 (n_10599, wc427, n_9420);
  not gc427 (wc427, n_10123);
  or g28214 (n_10586, wc428, n_9420);
  not gc428 (wc428, n_10195);
  or g28215 (n_10550, wc429, n_9420);
  not gc429 (wc429, n_10138);
  or g28216 (n_10568, wc430, n_9420);
  not gc430 (wc430, n_10156);
  or g28217 (n_9426, n_9411, wc431);
  not gc431 (wc431, n_9425);
  or g28218 (n_10585, wc432, n_9425);
  not gc432 (wc432, n_10196);
  or g28219 (n_10549, wc433, n_9425);
  not gc433 (wc433, n_10139);
  or g28220 (n_10567, wc434, n_9425);
  not gc434 (wc434, n_10157);
  or g28221 (n_10598, n_12840, n_9426);
  or g28222 (n_9428, wc435, n_10601);
  not gc435 (wc435, n_10600);
  or g28223 (n_9463, n_9346, wc436);
  not gc436 (wc436, n_9434);
  or g28224 (n_10607, wc437, n_9434);
  not gc437 (wc437, n_9346);
  or g28225 (n_10610, n_9357, wc438);
  not gc438 (wc438, n_9441);
  or g28226 (n_9900, wc439, n_9441);
  not gc439 (wc439, n_9357);
  or g28227 (n_9462, wc440, n_9447);
  not gc440 (wc440, n_9349);
  or g28228 (n_9944, n_9349, wc441);
  not gc441 (wc441, n_9447);
  or g28230 (n_12810, wc442, n_9429);
  not gc442 (wc442, n_9448);
  or g28232 (n_9470, n_9383, wc443);
  not gc443 (wc443, n_10685);
  or g28233 (n_9471, wc444, n_9449);
  not gc444 (wc444, n_9470);
  or g28234 (n_9461, n_9458, wc445);
  not gc445 (wc445, n_9449);
  or g28235 (n_9459, n_9419, wc446);
  not gc446 (wc446, n_9458);
  or g28236 (n_10715, n_12810, n_9471);
  or g28237 (n_9981, n_9459, wc447);
  not gc447 (wc447, n_9802);
  or g28238 (n_9516, n_9379, wc448);
  not gc448 (wc448, n_10706);
  or g28239 (n_9472, wc449, n_10718);
  not gc449 (wc449, n_10717);
  or g28240 (n_9869, n_9355, wc450);
  not gc450 (wc450, n_9499);
  or g28241 (n_10835, n_9352, wc451);
  not gc451 (wc451, n_9476);
  or g28242 (n_9931, wc452, n_9476);
  not gc452 (wc452, n_9352);
  or g28243 (n_10832, n_9349, wc453);
  not gc453 (wc453, n_9493);
  or g28244 (n_9936, wc454, n_9493);
  not gc454 (wc454, n_9349);
  or g28245 (n_10838, n_9346, wc455);
  not gc455 (wc455, n_9480);
  or g28246 (n_9965, wc456, n_9480);
  not gc456 (wc456, n_9346);
  or g28247 (n_10841, n_9357, wc457);
  not gc457 (wc457, n_9487);
  or g28248 (n_10002, wc458, n_9487);
  not gc458 (wc458, n_9357);
  or g28249 (n_10829, wc459, n_9499);
  not gc459 (wc459, n_9355);
  or g28250 (n_12194, wc460, n_9522);
  not gc460 (wc460, n_9869);
  or g28251 (n_10902, wc461, n_9500);
  not gc461 (wc461, n_10072);
  or g28252 (n_10906, wc462, n_10905);
  not gc462 (wc462, n_10904);
  or g28253 (n_11026, wc463, n_9524);
  not gc463 (wc463, n_10184);
  or g28254 (n_10990, wc464, n_9524);
  not gc464 (wc464, n_10169);
  or g28255 (n_10972, wc465, n_9524);
  not gc465 (wc465, n_10163);
  or g28256 (n_11044, wc466, n_9524);
  not gc466 (wc466, n_10202);
  or g28257 (n_11008, wc467, n_9524);
  not gc467 (wc467, n_10178);
  or g28258 (n_10954, wc468, n_9524);
  not gc468 (wc468, n_10154);
  or g28259 (n_10936, wc469, n_9524);
  not gc469 (wc469, n_10133);
  or g28260 (n_10146, wc470, n_12260);
  not gc470 (wc470, n_12259);
  or g28261 (n_9525, wc471, n_9501);
  not gc471 (wc471, n_9524);
  or g28262 (n_9512, wc472, n_9846);
  not gc472 (wc472, n_10146);
  or g28263 (n_10919, wc473, n_9514);
  not gc473 (wc473, n_10119);
  or g28264 (n_11025, wc474, n_9514);
  not gc474 (wc474, n_10185);
  or g28265 (n_10989, wc475, n_9514);
  not gc475 (wc475, n_10170);
  or g28266 (n_10971, wc476, n_9514);
  not gc476 (wc476, n_10164);
  or g28267 (n_11043, wc477, n_9514);
  not gc477 (wc477, n_10203);
  or g28268 (n_11007, wc478, n_9514);
  not gc478 (wc478, n_10179);
  or g28269 (n_10953, wc479, n_9514);
  not gc479 (wc479, n_10155);
  or g28270 (n_10935, wc480, n_9514);
  not gc480 (wc480, n_10134);
  or g28271 (n_9527, wc481, n_10922);
  not gc481 (wc481, n_10921);
  or g28272 (n_11060, wc482, n_9533);
  not gc482 (wc482, n_9381);
  or g28273 (n_11057, n_9355, wc483);
  not gc483 (wc483, n_9567);
  or g28274 (n_9954, wc484, n_9567);
  not gc484 (wc484, n_9355);
  or g28275 (n_11063, n_9352, wc485);
  not gc485 (wc485, n_9544);
  or g28276 (n_9910, wc486, n_9544);
  not gc486 (wc486, n_9352);
  or g28277 (n_11054, n_9349, wc487);
  not gc487 (wc487, n_9561);
  or g28278 (n_9897, wc488, n_9561);
  not gc488 (wc488, n_9349);
  or g28279 (n_11066, n_9346, wc489);
  not gc489 (wc489, n_9548);
  or g28280 (n_9907, wc490, n_9548);
  not gc490 (wc490, n_9346);
  or g28281 (n_11069, n_9357, wc491);
  not gc491 (wc491, n_9555);
  or g28282 (n_9961, wc492, n_9555);
  not gc492 (wc492, n_9357);
  or g28283 (n_9585, wc493, n_9538);
  not gc493 (wc493, n_9382);
  or g28284 (n_11051, n_9382, wc494);
  not gc494 (wc494, n_9538);
  or g28285 (n_9586, wc495, n_9381);
  not gc495 (wc495, n_9533);
  or g28286 (n_12328, wc496, n_9596);
  not gc496 (wc496, n_11125);
  or g28287 (n_12329, n_12328, wc497);
  not gc497 (wc497, n_9839);
  or g28288 (n_10204, n_12329, wc498);
  not gc498 (wc498, n_9585);
  or g28289 (n_9866, wc499, n_12344);
  not gc499 (wc499, n_12343);
  or g28290 (n_11206, wc500, n_9597);
  not gc500 (wc500, n_10130);
  or g28291 (n_11224, wc501, n_9597);
  not gc501 (wc501, n_10136);
  or g28292 (n_11242, wc502, n_9597);
  not gc502 (wc502, n_10142);
  or g28293 (n_11347, wc503, n_9597);
  not gc503 (wc503, n_10199);
  or g28294 (n_11293, wc504, n_9597);
  not gc504 (wc504, n_10166);
  or g28295 (n_11311, wc505, n_9597);
  not gc505 (wc505, n_10172);
  or g28296 (n_11329, wc506, n_9597);
  not gc506 (wc506, n_10175);
  or g28297 (n_11275, wc507, n_9597);
  not gc507 (wc507, n_10151);
  or g28298 (n_11188, wc508, n_9597);
  not gc508 (wc508, n_10127);
  or g28299 (n_9583, n_9513, wc509);
  not gc509 (wc509, n_9582);
  or g28300 (n_9598, wc510, n_9570);
  not gc510 (wc510, n_9597);
  or g28301 (n_9584, n_9582, wc511);
  not gc511 (wc511, n_9570);
  or g28302 (n_9600, wc512, n_11261);
  not gc512 (wc512, n_11260);
  or g28303 (n_9667, n_9377, wc513);
  not gc513 (wc513, n_9604);
  or g28304 (n_9668, wc514, n_9608);
  not gc514 (wc514, n_9382);
  or g28305 (n_9678, n_9381, wc515);
  not gc515 (wc515, n_9612);
  or g28306 (n_9669, wc516, n_9612);
  not gc516 (wc516, n_9381);
  or g28307 (n_11360, n_9355, wc517);
  not gc517 (wc517, n_9639);
  or g28308 (n_9983, wc518, n_9639);
  not gc518 (wc518, n_9355);
  or g28309 (n_11363, n_9352, wc519);
  not gc519 (wc519, n_9616);
  or g28310 (n_9979, wc520, n_9616);
  not gc520 (wc520, n_9352);
  or g28311 (n_11366, n_9349, wc521);
  not gc521 (wc521, n_9633);
  or g28312 (n_9985, wc522, n_9633);
  not gc522 (wc522, n_9349);
  or g28313 (n_11369, n_9346, wc523);
  not gc523 (wc523, n_9620);
  or g28314 (n_9902, wc524, n_9620);
  not gc524 (wc524, n_9346);
  or g28315 (n_11357, n_9357, wc525);
  not gc525 (wc525, n_9627);
  or g28316 (n_9964, wc526, n_9627);
  not gc526 (wc526, n_9357);
  or g28317 (n_9908, n_9382, wc527);
  not gc527 (wc527, n_9608);
  or g28318 (n_9683, wc528, n_9648);
  not gc528 (wc528, n_9378);
  or g28319 (n_9652, wc529, n_9604);
  not gc529 (wc529, n_9377);
  or g28320 (n_9881, n_9378, wc530);
  not gc530 (wc530, n_9648);
  or g28321 (n_10071, b12, wc531);
  not gc531 (wc531, n_11354);
  or g28322 (n_9838, wc532, n_9679);
  not gc532 (wc532, n_9652);
  or g28323 (n_11447, wc533, n_9677);
  not gc533 (wc533, n_9668);
  or g28324 (n_9684, n_11447, wc534);
  not gc534 (wc534, n_9652);
  or g28325 (n_11459, wc535, n_11457);
  not gc535 (wc535, n_9686);
  or g28326 (n_11644, wc536, n_9687);
  not gc536 (wc536, n_10102);
  or g28327 (n_9688, wc537, n_9650);
  not gc537 (wc537, n_9687);
  or g28328 (n_11536, wc538, n_9687);
  not gc538 (wc538, n_10081);
  or g28329 (n_11590, wc539, n_9687);
  not gc539 (wc539, n_10090);
  or g28330 (n_11626, wc540, n_9687);
  not gc540 (wc540, n_10099);
  or g28331 (n_11662, wc541, n_9687);
  not gc541 (wc541, n_10105);
  or g28332 (n_11716, wc542, n_9687);
  not gc542 (wc542, n_10114);
  or g28333 (n_11698, wc543, n_9687);
  not gc543 (wc543, n_10111);
  or g28334 (n_11680, wc544, n_9687);
  not gc544 (wc544, n_10108);
  or g28335 (n_11608, wc545, n_9687);
  not gc545 (wc545, n_10096);
  or g28336 (n_11572, wc546, n_9687);
  not gc546 (wc546, n_10087);
  or g28337 (n_11554, wc547, n_9687);
  not gc547 (wc547, n_10084);
  or g28338 (n_9695, n_9583, wc548);
  not gc548 (wc548, n_9665);
  or g28339 (n_11643, wc549, n_9666);
  not gc549 (wc549, n_10103);
  or g28340 (n_11535, wc550, n_9666);
  not gc550 (wc550, n_10082);
  or g28341 (n_11589, wc551, n_9666);
  not gc551 (wc551, n_10091);
  or g28342 (n_11625, wc552, n_9666);
  not gc552 (wc552, n_10100);
  or g28343 (n_11661, wc553, n_9666);
  not gc553 (wc553, n_10106);
  or g28344 (n_11519, wc554, n_9666);
  not gc554 (wc554, n_10077);
  or g28345 (n_11715, wc555, n_9666);
  not gc555 (wc555, n_10115);
  or g28346 (n_11697, wc556, n_9666);
  not gc556 (wc556, n_10112);
  or g28347 (n_11679, wc557, n_9666);
  not gc557 (wc557, n_10109);
  or g28348 (n_11607, wc558, n_9666);
  not gc558 (wc558, n_10097);
  or g28349 (n_11571, wc559, n_9666);
  not gc559 (wc559, n_10088);
  or g28350 (n_11553, wc560, n_9666);
  not gc560 (wc560, n_10085);
  or g28351 (n_9698, wc561, n_11522);
  not gc561 (wc561, n_11521);
  or g28352 (n_9853, wc562, n_9694);
  not gc562 (wc562, n_9372);
  or g28353 (n_10030, wc563, n_9739);
  not gc563 (wc563, n_9349);
  or g28354 (n_10040, wc564, n_9719);
  not gc564 (wc564, n_9382);
  or g28355 (n_10062, wc565, n_9705);
  not gc565 (wc565, n_9378);
  or g28356 (n_10063, wc566, n_9708);
  not gc566 (wc566, n_9377);
  or g28357 (n_10064, wc567, n_9725);
  not gc567 (wc567, n_9352);
  or g28358 (n_10065, wc568, n_9729);
  not gc568 (wc568, n_9355);
  or g28359 (n_11764, n_9372, wc569);
  not gc569 (wc569, n_9694);
  or g28360 (n_11896, wc570, n_9705);
  not gc570 (wc570, n_9377);
  or g28361 (n_11753, n_9382, wc571);
  not gc571 (wc571, n_9715);
  or g28362 (n_11875, wc572, n_9729);
  not gc572 (wc572, n_9352);
  or g28363 (n_11756, n_9349, wc573);
  not gc573 (wc573, n_9735);
  or g28364 (n_12435, wc574, n_9748);
  not gc574 (wc574, n_9357);
  or g28365 (n_11866, wc575, n_9689);
  not gc575 (wc575, n_9371);
  or g28366 (n_11774, n_9328, wc576);
  not gc576 (wc576, n_9715);
  or g28367 (n_11787, n_9326, wc577);
  not gc577 (wc577, n_9735);
  or g28368 (n_11763, wc578, n_9371);
  not gc578 (wc578, n_9853);
  or g28369 (n_12434, wc579, n_9745);
  not gc579 (wc579, n_9400);
  or g28370 (n_11900, n_9400, wc580);
  not gc580 (wc580, n_9745);
  or g28371 (n_11926, n_9689, wc581);
  not gc581 (wc581, n_9843);
  or g28372 (n_11948, n_9338, wc582);
  not gc582 (wc582, n_9745);
  or g28373 (n_11765, n_11763, wc583);
  not gc583 (wc583, n_9689);
  or g28374 (n_11990, wc584, n_9767);
  not gc584 (wc584, n_9735);
  or g28375 (n_11996, wc585, n_9760);
  not gc585 (wc585, n_9715);
  or g28376 (n_9740, n_11834, wc586);
  not gc586 (wc586, n_9731);
  or g28377 (n_11968, wc587, n_9815);
  not gc587 (wc587, n_10023);
  or g28378 (n_11977, wc588, n_9812);
  not gc588 (wc588, n_10024);
  or g28379 (n_12437, wc589, n_12436);
  not gc589 (wc589, n_12435);
  or g28380 (n_10037, wc590, n_11813);
  not gc590 (wc590, n_11812);
  or g28381 (n_11916, n_9740, wc591);
  not gc591 (wc591, n_9735);
  or g28382 (n_10032, wc592, n_11777);
  not gc592 (wc592, n_11776);
  or g28383 (n_10033, wc593, n_11789);
  not gc593 (wc593, n_11788);
  or g28384 (n_9769, n_12437, wc594);
  not gc594 (wc594, n_11857);
  or g28385 (n_9720, wc595, n_9711);
  not gc595 (wc595, n_10037);
  or g28386 (n_10009, n_11741, wc596);
  not gc596 (wc596, n_9359);
  or g28387 (n_9780, wc597, n_9775);
  not gc597 (wc597, n_10032);
  or g28388 (n_9785, wc598, n_9782);
  not gc598 (wc598, n_10033);
  or g28389 (n_9762, wc599, n_9761);
  not gc599 (wc599, n_10021);
  or g28390 (n_9772, wc600, n_9771);
  not gc600 (wc600, n_10011);
  or g28391 (n_9770, wc601, n_11960);
  not gc601 (wc601, n_11959);
  or g28392 (n_9721, n_9710, wc602);
  not gc602 (wc602, n_11993);
  or g28393 (n_9742, wc603, n_9741);
  not gc603 (wc603, n_10034);
  or g28394 (n_12017, wc604, n_12016);
  not gc604 (wc604, n_9770);
  or g28395 (n_9787, n_9786, wc605);
  not gc605 (wc605, n_12011);
  or g28396 (n_12025, wc606, n_12024);
  not gc606 (wc606, n_9787);
  or g28397 (n_10042, n_9762, wc607);
  not gc607 (wc607, n_12038);
  or g28398 (n_12062, wc608, n_9764);
  not gc608 (wc608, n_10042);
  or g28399 (n_12058, wc609, n_12057);
  not gc609 (wc609, n_12056);
  or g28400 (n_10045, n_9781, wc610);
  not gc610 (wc610, n_12026);
  or g28401 (n_12041, wc611, n_9777);
  not gc611 (wc611, n_10045);
  or g28402 (n_9751, b15, wc612);
  not gc612 (wc612, n_12071);
  and g28403 (o1, wc613, n_9335);
  not gc613 (wc613, n_9751);
endmodule

