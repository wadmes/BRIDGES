module test(a7, a6, a5, a4, a3, a2, a1, a0, b7, b6, b5, b4, b3, b2, b1,
     b0, o7, o6, o5, o4, o3, o2, o1, o0);
  input a7, a6, a5, a4, a3, a2, a1, a0, b7, b6, b5, b4, b3, b2, b1, b0;
  output o7, o6, o5, o4, o3, o2, o1, o0;
  wire a7, a6, a5, a4, a3, a2, a1, a0, b7, b6, b5, b4, b3, b2, b1, b0;
  wire o7, o6, o5, o4, o3, o2, o1, o0;
  wire anoymous_7_126_n_25, anoymous_7_126_n_26, anoymous_7_126_n_27, anoymous_7_126_n_28,
       anoymous_7_126_n_29, anoymous_7_126_n_30, anoymous_7_126_n_31, anoymous_7_126_n_40;
  wire anoymous_7_126_n_47, anoymous_7_126_n_48, anoymous_7_126_n_59, anoymous_7_126_n_61,
       anoymous_7_126_n_62, anoymous_7_126_n_64, anoymous_7_126_n_68, anoymous_7_126_n_69;
  wire anoymous_7_126_n_70, anoymous_7_126_n_71, anoymous_7_126_n_89, anoymous_7_126_n_90,
       anoymous_7_126_n_91, anoymous_7_126_n_93, anoymous_7_126_n_94, anoymous_7_126_n_97;
  wire anoymous_7_126_n_98, anoymous_7_126_n_99, anoymous_7_126_n_100,
       anoymous_7_126_n_101, anoymous_7_126_n_102, anoymous_7_126_n_127,
       anoymous_7_126_n_133, anoymous_7_126_n_152;
  wire anoymous_7_126_n_156, anoymous_7_126_n_162, anoymous_7_126_n_166,
       anoymous_7_126_n_167, anoymous_7_126_n_181, anoymous_7_126_n_193,
       anoymous_7_126_n_196, anoymous_7_126_n_200;
  wire anoymous_7_126_n_202, anoymous_7_126_n_316, anoymous_7_126_n_322,
       anoymous_7_126_n_340, anoymous_7_126_n_350, anoymous_7_126_n_368,
       anoymous_7_126_n_388, anoymous_7_126_n_495;
  wire anoymous_7_126_n_511, anoymous_7_126_n_524, anoymous_7_126_n_536,
       anoymous_7_126_n_537, anoymous_7_126_n_539, anoymous_7_126_n_540,
       anoymous_7_126_n_541, anoymous_7_126_n_559;
  wire anoymous_7_126_n_589, anoymous_7_126_n_604, anoymous_7_126_n_606,
       anoymous_7_126_n_607, anoymous_7_126_n_643, anoymous_7_126_n_658,
       anoymous_7_126_n_672, anoymous_7_126_n_673;
  wire anoymous_7_126_n_675, anoymous_7_126_n_676, anoymous_7_126_n_723,
       anoymous_7_126_n_729, anoymous_7_126_n_732, anoymous_7_126_n_734,
       anoymous_7_126_n_806, anoymous_7_126_n_809;
  wire anoymous_7_126_n_811, anoymous_7_126_n_821, anoymous_7_126_n_879,
       anoymous_7_126_n_885, n_46, n_1469, n_1820, n_1821;
  wire n_1835, n_1845, n_1848, n_1849, n_1850, n_1852, n_1855, n_1856;
  wire n_1857, n_1858, n_1861, n_1862, n_1863, n_1864, n_1865, n_1866;
  wire n_1868, n_1870, n_1871, n_1873, n_1874, n_1876, n_1879, n_1880;
  wire n_1883, n_1885, n_1887, n_1889, n_1892, n_1893, n_1895, n_1896;
  wire n_1897, n_1898, n_1905, n_1911, n_1916, n_1917, n_1919, n_1920;
  wire n_1921, n_1922, n_1923, n_1925, n_1926, n_1927, n_1928, n_1929;
  wire n_1930, n_1931, n_1932, n_1934, n_1935, n_1936, n_1938, n_1939;
  wire n_1940, n_1941, n_1942, n_1943, n_1944, n_1945, n_1946, n_1947;
  wire n_1948, n_1949, n_1950, n_1951, n_1952, n_1953, n_1954, n_1955;
  wire n_1956, n_1958, n_1959, n_1960, n_1961, n_1962, n_1964, n_1965;
  wire n_1967, n_1968, n_1972, n_1975, n_1978, n_1981, n_1984, n_1987;
  wire n_1992, n_1993, n_2002, n_2003, n_2010, n_2011, n_2016, n_2017;
  wire n_2020, n_2023, n_2026, n_2037, n_2039, n_2040, n_2041, n_2058;
  wire n_2059, n_2060, n_2061, n_2062, n_2063, n_2064, n_2073, n_2074;
  wire n_2089, n_2090, n_2091, n_2092, n_2093, n_2094, n_2095, n_2108;
  wire n_2109, n_2110, n_2111, n_2112, n_2113, n_2122, n_2123, n_2124;
  wire n_2125, n_2128, n_2131, n_2134, n_2137, n_2140, n_2143, n_2146;
  wire n_2149, n_2156, n_2158, n_2169, n_2170, n_2171, n_2172, n_2178;
  wire n_2179, n_2192, n_2193, n_2194, n_2195, n_2196, n_2197, n_2210;
  wire n_2211, n_2212, n_2213, n_2214, n_2215, n_2228, n_2229, n_2230;
  wire n_2231, n_2232, n_2233, n_2246, n_2247, n_2248, n_2249, n_2250;
  wire n_2251, n_2260, n_2261, n_2262, n_2263, n_2270, n_2271, n_2272;
  wire n_2283, n_2284, n_2285, n_2286, n_2287, n_2294, n_2295, n_2296;
  wire n_2299, n_2302, n_2309, n_2310, n_2311, n_2320, n_2321, n_2322;
  wire n_2323, n_2332, n_2333, n_2334, n_2335, n_2340, n_2341, n_2352;
  wire n_2353, n_2354, n_2355, n_2356, n_2361, n_2362, n_2380, n_2381;
  wire n_2382, n_2383, n_2384, n_2385, n_2386, n_2391, n_2392, n_2397;
  wire n_2398, n_2401, n_2404, n_2407, n_2412, n_2413, n_2416, n_2423;
  wire n_2424, n_2425, n_2436, n_2437, n_2438, n_2439, n_2440, n_2447;
  wire n_2448, n_2449, n_2452, n_2455, n_2458, n_2461, n_2464, n_2467;
  wire n_2476, n_2477, n_2478, n_2479, n_2482, n_2495, n_2496, n_2497;
  wire n_2498, n_2499, n_2500, n_2587, n_2589, n_2598, n_2599, n_2602;
  wire n_2603, n_2604, n_2606, n_2607, n_2608, n_2609, n_2610, n_2611;
  wire n_2612, n_2613, n_2614, n_2615, n_2616, n_2617, n_2618, n_2619;
  wire n_2622, n_2623, n_2625, n_2629, n_2630, n_2631, n_2632, n_2634;
  wire n_2635, n_2636, n_2638, n_2639, n_2640, n_2641, n_2642, n_2643;
  wire n_2644, n_2645, n_2646, n_2647, n_2648, n_2649, n_2650, n_2651;
  wire n_2652, n_2653;
  or g2878 (anoymous_7_126_n_340, wc, a4);
  not gc (wc, b0);
  or g2884 (anoymous_7_126_n_495, wc0, a2);
  not gc0 (wc0, b0);
  or g3722 (n_1820, b3, wc1);
  not gc1 (wc1, anoymous_7_126_n_70);
  or g3974 (n_1855, b5, b6);
  or g3975 (n_1835, n_1855, b7);
  nand g3984 (n_1857, b3, b2);
  nand g3990 (n_1858, b4, b3);
  nand g3999 (n_1861, b5, b4);
  or g4025 (n_1868, anoymous_7_126_n_25, wc2);
  not gc2 (wc2, a5);
  nand g4031 (n_1870, b1, b0);
  or g4050 (n_1876, anoymous_7_126_n_495, a3);
  or g4102 (n_1892, wc3, a5);
  not gc3 (wc3, b1);
  or g4103 (n_1885, b1, wc4);
  not gc4 (wc4, a7);
  or g4104 (n_1856, wc5, a6);
  not gc5 (wc5, b0);
  or g4134 (n_1895, wc6, anoymous_7_126_n_69);
  not gc6 (wc6, b3);
  or g4135 (n_1866, wc7, anoymous_7_126_n_70);
  not gc7 (wc7, b4);
  or g4136 (n_1887, wc8, anoymous_7_126_n_69);
  not gc8 (wc8, b2);
  or g4137 (n_1896, wc9, anoymous_7_126_n_68);
  not gc9 (wc9, b2);
  or g4141 (n_1880, wc10, anoymous_7_126_n_68);
  not gc10 (wc10, b1);
  or g4163 (n_1850, wc11, anoymous_7_126_n_100);
  not gc11 (wc11, b5);
  or g4166 (n_1873, wc12, anoymous_7_126_n_98);
  not gc12 (wc12, b3);
  nand g4383 (n_1911, n_1821, n_1865);
  nand g4416 (n_1925, b0, n_1862);
  nand g4419 (n_1926, b0, n_1863);
  or g4422 (n_1927, anoymous_7_126_n_31, anoymous_7_126_n_30);
  or g4535 (n_1941, anoymous_7_126_n_101, wc13);
  not gc13 (wc13, b5);
  or g4541 (n_1944, anoymous_7_126_n_101, wc14);
  not gc14 (wc14, b6);
  or g4549 (n_1948, anoymous_7_126_n_28, wc15);
  not gc15 (wc15, anoymous_7_126_n_70);
  nand g4581 (n_1964, n_1469, b0);
  nand g5031 (n_1930, anoymous_7_126_n_133, n_2404);
  nand g5032 (n_2404, anoymous_7_126_n_322, n_1883);
  or g5033 (n_1883, n_2499, n_2500);
  nand g5034 (n_2499, n_2495, n_2496);
  or g5035 (n_2496, wc16, anoymous_7_126_n_885);
  not gc16 (wc16, n_1939);
  nand g5038 (n_1939, n_2397, n_2398);
  nand g5039 (anoymous_7_126_n_133, n_1938, anoymous_7_126_n_127);
  nand g5040 (n_2397, n_1849, n_1916);
  or g5042 (n_1938, n_2385, n_2386);
  or g5043 (n_2401, wc17, anoymous_7_126_n_821);
  not gc17 (wc17, n_1942);
  nand g5044 (n_1916, n_2361, n_2362);
  or g5046 (n_1942, n_1917, n_2392);
  nand g5048 (n_2362, n_1936, anoymous_7_126_n_99);
  nand g5050 (anoymous_7_126_n_809, n_2322, n_2323);
  nand g5051 (n_2380, n_1923, anoymous_7_126_n_734);
  nand g5052 (anoymous_7_126_n_732, n_2310, n_2311);
  or g5053 (n_1936, n_2356, wc18);
  not gc18 (wc18, anoymous_7_126_n_28);
  or g5054 (n_2361, wc19, anoymous_7_126_n_28);
  not gc19 (wc19, n_2356);
  nand g5055 (n_2392, anoymous_7_126_n_811, n_2391);
  nand g5056 (n_1923, n_1898, n_2482);
  or g5057 (n_2356, n_2355, wc20);
  not gc20 (wc20, anoymous_7_126_n_879);
  nand g5058 (anoymous_7_126_n_811, n_2340, n_2341);
  or g5060 (n_2322, n_2320, b3);
  or g5061 (n_2310, n_1898, wc21);
  not gc21 (wc21, anoymous_7_126_n_99);
  or g5062 (n_2311, n_2309, b5);
  or g5063 (n_2482, n_2299, wc22);
  not gc22 (wc22, anoymous_7_126_n_99);
  or g5064 (n_2323, n_2321, b4);
  nand g5065 (n_2355, n_2353, n_2354);
  or g5066 (n_1898, n_2299, b4);
  nand g5067 (n_2341, n_1932, anoymous_7_126_n_98);
  or g5070 (n_1935, n_2272, wc23);
  not gc23 (wc23, n_1905);
  nand g5071 (n_2335, anoymous_7_126_n_723, n_2333);
  or g5072 (n_1917, anoymous_7_126_n_806, wc24);
  not gc24 (wc24, n_2302);
  nand g5073 (n_2272, n_2270, n_2271);
  or g5075 (n_1932, n_2296, wc25);
  not gc25 (wc25, b2);
  or g5076 (n_2299, wc26, anoymous_7_126_n_729);
  not gc26 (wc26, n_1850);
  or g5078 (n_2309, anoymous_7_126_n_729, wc27);
  not gc27 (wc27, anoymous_7_126_n_100);
  or g5079 (n_2354, n_2352, wc28);
  not gc28 (wc28, anoymous_7_126_n_97);
  or g5080 (n_2340, wc29, b2);
  not gc29 (wc29, n_2296);
  or g5081 (n_2334, n_2332, b2);
  or g5082 (n_2321, anoymous_7_126_n_806, wc30);
  not gc30 (wc30, anoymous_7_126_n_100);
  nand g5083 (n_2332, n_1873, anoymous_7_126_n_97);
  or g5084 (n_2383, n_1852, b6);
  or g5085 (n_2495, n_1852, anoymous_7_126_n_30);
  nand g5086 (anoymous_7_126_n_729, n_1944, n_1943);
  or g5087 (n_2352, anoymous_7_126_n_26, wc31);
  not gc31 (wc31, n_1871);
  nand g5088 (n_2271, n_1852, b6);
  nand g5089 (n_2500, n_2497, n_2498);
  nand g5090 (n_2478, n_2476, n_2477);
  nand g5091 (n_2296, n_2294, n_2295);
  nand g5092 (n_2385, n_2381, n_2382);
  or g5093 (n_2287, wc32, n_2286);
  not gc32 (wc32, n_2285);
  nand g5094 (anoymous_7_126_n_806, n_1941, n_1940);
  nand g5095 (anoymous_7_126_n_885, n_1929, n_1928);
  or g5096 (n_2302, anoymous_7_126_n_100, wc33);
  not gc33 (wc33, b4);
  or g5097 (n_2285, anoymous_7_126_n_97, wc34);
  not gc34 (wc34, b2);
  or g5098 (n_2333, wc35, b3);
  not gc35 (wc35, anoymous_7_126_n_98);
  or g5099 (n_2391, anoymous_7_126_n_99, wc36);
  not gc36 (wc36, b3);
  or g5100 (n_2498, n_1927, wc37);
  not gc37 (wc37, anoymous_7_126_n_101);
  nand g5105 (n_2294, n_1931, anoymous_7_126_n_97);
  or g5108 (anoymous_7_126_n_100, n_2250, n_2251);
  or g5109 (anoymous_7_126_n_99, n_2214, n_2215);
  nand g5110 (n_2598, n_1925, a2);
  or g5111 (n_2599, n_1925, a2);
  nand g5112 (anoymous_7_126_n_97, n_2598, n_2599);
  or g5113 (anoymous_7_126_n_98, n_2232, n_2233);
  or g5114 (anoymous_7_126_n_101, n_2263, wc38);
  not gc38 (wc38, n_2262);
  nand g5117 (n_2233, n_2230, n_2231);
  nand g5118 (n_2263, n_2260, n_2261);
  nand g5119 (n_2251, n_2248, n_2249);
  nand g5120 (n_2232, n_2228, n_2229);
  nand g5121 (n_2214, n_2210, n_2211);
  nand g5122 (n_2250, n_2246, n_2247);
  nand g5123 (n_2215, n_2212, n_2213);
  or g5124 (n_2230, wc39, anoymous_7_126_n_91);
  not gc39 (wc39, n_1950);
  nand g5125 (n_2270, n_1934, b5);
  or g5126 (n_2261, wc40, anoymous_7_126_n_91);
  not gc40 (wc40, n_1962);
  or g5128 (n_2247, wc41, anoymous_7_126_n_94);
  not gc41 (wc41, n_1960);
  or g5129 (n_2248, wc42, anoymous_7_126_n_91);
  not gc42 (wc42, n_1959);
  or g5130 (n_2212, wc43, anoymous_7_126_n_91);
  not gc43 (wc43, n_1953);
  or g5131 (n_2211, wc44, anoymous_7_126_n_94);
  not gc44 (wc44, n_1954);
  or g5132 (n_2229, wc45, anoymous_7_126_n_94);
  not gc45 (wc45, n_1951);
  nand g5133 (n_1862, anoymous_7_126_n_91, anoymous_7_126_n_93);
  nand g5134 (n_1940, anoymous_7_126_n_102, b6);
  or g5135 (n_1934, anoymous_7_126_n_102, b6);
  or g5136 (n_2497, anoymous_7_126_n_31, anoymous_7_126_n_102);
  nand g5139 (n_1928, anoymous_7_126_n_31, anoymous_7_126_n_102);
  or g5140 (n_2382, anoymous_7_126_n_102, b7);
  nand g5141 (n_1943, anoymous_7_126_n_102, b7);
  nand g5145 (n_2231, anoymous_7_126_n_89, a3);
  nand g5146 (n_2262, anoymous_7_126_n_89, anoymous_7_126_n_70);
  nand g5147 (n_2213, anoymous_7_126_n_68, anoymous_7_126_n_89);
  or g5148 (anoymous_7_126_n_90, n_1835, n_2197);
  nand g5149 (n_2249, anoymous_7_126_n_89, anoymous_7_126_n_69);
  or g5151 (anoymous_7_126_n_89, wc46, anoymous_7_126_n_166);
  not gc46 (wc46, n_1958);
  nand g5155 (n_1958, n_2178, n_2179);
  nand g5156 (n_2196, n_2193, n_2194);
  or g5158 (anoymous_7_126_n_93, n_1927, n_2172);
  nand g5159 (n_2193, anoymous_7_126_n_71, n_1945);
  or g5160 (n_2179, wc47, anoymous_7_126_n_71);
  not gc47 (wc47, n_1956);
  nand g5161 (n_2172, n_2170, n_2171);
  or g5162 (n_1956, n_2158, wc48);
  not gc48 (wc48, b5);
  or g5163 (n_2178, wc49, b5);
  not gc49 (wc49, n_2158);
  or g5164 (n_1945, n_2467, b4);
  nand g5165 (n_2158, n_2156, n_2134);
  or g5166 (n_2195, n_2192, wc50);
  not gc50 (wc50, b4);
  nand g5167 (n_2467, n_2192, n_2128);
  or g5169 (n_2192, wc51, anoymous_7_126_n_589);
  not gc51 (wc51, n_1820);
  nand g5170 (n_2156, n_1866, anoymous_7_126_n_524);
  nand g5171 (n_2602, anoymous_7_126_n_541, anoymous_7_126_n_524);
  or g5172 (n_2603, anoymous_7_126_n_541, anoymous_7_126_n_524);
  nand g5173 (n_1962, n_2602, n_2603);
  nand g5178 (anoymous_7_126_n_524, n_2140, n_2455);
  nand g5179 (n_2449, n_2447, n_2448);
  nand g5180 (anoymous_7_126_n_589, n_2137, n_2452);
  nand g5182 (n_2606, anoymous_7_126_n_676, anoymous_7_126_n_675);
  or g5183 (n_2607, anoymous_7_126_n_676, anoymous_7_126_n_675);
  nand g5184 (n_1961, n_2606, n_2607);
  nand g5185 (n_2608, anoymous_7_126_n_540, anoymous_7_126_n_539);
  or g5186 (n_2609, anoymous_7_126_n_540, anoymous_7_126_n_539);
  nand g5187 (n_1959, n_2608, n_2609);
  nand g5188 (n_2455, n_1895, anoymous_7_126_n_539);
  nand g5189 (n_2610, anoymous_7_126_n_607, anoymous_7_126_n_606);
  or g5190 (n_2611, anoymous_7_126_n_607, anoymous_7_126_n_606);
  nand g5191 (n_1960, n_2610, n_2611);
  nand g5192 (n_2452, n_1887, anoymous_7_126_n_606);
  nand g5193 (anoymous_7_126_n_606, n_2149, n_2464);
  nand g5194 (n_2612, anoymous_7_126_n_511, anoymous_7_126_n_537);
  or g5195 (n_2613, anoymous_7_126_n_511, anoymous_7_126_n_537);
  nand g5196 (n_1953, n_2612, n_2613);
  nand g5197 (anoymous_7_126_n_539, n_2143, n_2458);
  or g5198 (n_2614, anoymous_7_126_n_559, anoymous_7_126_n_604);
  nand g5199 (n_2615, anoymous_7_126_n_559, anoymous_7_126_n_604);
  nand g5200 (n_1954, n_2614, n_2615);
  nand g5201 (n_2616, anoymous_7_126_n_643, anoymous_7_126_n_673);
  or g5202 (n_2617, anoymous_7_126_n_643, anoymous_7_126_n_673);
  nand g5203 (n_1955, n_2616, n_2617);
  nand g5204 (anoymous_7_126_n_675, n_2146, n_2461);
  nand g5205 (anoymous_7_126_n_673, n_1893, n_2146);
  nand g5206 (n_2169, n_1949, n_1948);
  nand g5207 (anoymous_7_126_n_676, n_1889, n_2131);
  nand g5208 (anoymous_7_126_n_604, n_1880, n_2149);
  nand g5209 (n_2464, anoymous_7_126_n_559, n_1880);
  nand g5210 (anoymous_7_126_n_540, n_1895, n_2140);
  nand g5212 (n_2461, anoymous_7_126_n_643, n_1893);
  nand g5213 (anoymous_7_126_n_537, n_1896, n_2143);
  nand g5214 (anoymous_7_126_n_607, n_1887, n_2137);
  nand g5215 (n_2458, anoymous_7_126_n_511, n_1896);
  nand g5216 (anoymous_7_126_n_541, n_1866, n_2134);
  or g5217 (n_2447, wc52, anoymous_7_126_n_70);
  not gc52 (wc52, anoymous_7_126_n_28);
  or g5218 (n_2134, wc53, b4);
  not gc53 (wc53, anoymous_7_126_n_70);
  or g5219 (n_2137, wc54, b2);
  not gc54 (wc54, anoymous_7_126_n_69);
  or g5220 (n_2140, wc55, b3);
  not gc55 (wc55, anoymous_7_126_n_69);
  or g5222 (n_2143, wc56, b2);
  not gc56 (wc56, anoymous_7_126_n_68);
  or g5224 (n_2149, wc57, b1);
  not gc57 (wc57, anoymous_7_126_n_68);
  or g5225 (n_2128, anoymous_7_126_n_70, wc58);
  not gc58 (wc58, b3);
  or g5226 (n_2194, n_1858, anoymous_7_126_n_70);
  nand g5227 (n_2618, n_1926, a4);
  or g5228 (n_2619, n_1926, a4);
  nand g5229 (anoymous_7_126_n_68, n_2618, n_2619);
  or g5230 (anoymous_7_126_n_69, n_2112, n_2113);
  nand g5232 (n_2113, n_2110, n_2111);
  nand g5235 (n_2125, n_2122, n_2123);
  nand g5236 (n_2170, anoymous_7_126_n_71, anoymous_7_126_n_29);
  nand g5237 (n_1863, anoymous_7_126_n_62, anoymous_7_126_n_64);
  or g5238 (n_2123, wc59, anoymous_7_126_n_62);
  not gc59 (wc59, n_1965);
  or g5239 (n_2110, wc60, anoymous_7_126_n_62);
  not gc60 (wc60, n_1967);
  or g5240 (n_1949, anoymous_7_126_n_71, anoymous_7_126_n_29);
  nand g5241 (n_2112, n_2108, n_2109);
  nand g5243 (n_2111, anoymous_7_126_n_59, a5);
  or g5247 (n_2109, wc61, n_1879);
  not gc61 (wc61, n_1968);
  or g5248 (anoymous_7_126_n_59, n_1845, n_2440);
  nand g5253 (n_2439, n_2436, n_2437);
  or g5254 (anoymous_7_126_n_61, n_2095, anoymous_7_126_n_152);
  or g5256 (n_2095, n_1835, n_2094);
  nand g5258 (n_2437, n_1947, anoymous_7_126_n_48);
  or g5259 (n_1947, n_2074, b3);
  or g5260 (n_2094, wc62, n_2093);
  not gc62 (wc62, n_2092);
  or g5261 (anoymous_7_126_n_64, n_2064, anoymous_7_126_n_316);
  nand g5262 (n_2622, anoymous_7_126_n_350, n_1911);
  or g5263 (n_2623, anoymous_7_126_n_350, n_1911);
  nand g5264 (n_1965, n_2622, n_2623);
  or g5265 (n_2436, n_2073, wc63);
  not gc63 (wc63, b3);
  nand g5269 (n_2074, n_1865, n_2073);
  or g5270 (n_2092, n_2089, anoymous_7_126_n_388);
  or g5271 (n_2064, n_2062, n_2063);
  nand g5272 (n_2089, n_1921, n_1874);
  or g5273 (n_2073, wc64, anoymous_7_126_n_350);
  not gc64 (wc64, n_1821);
  nand g5274 (n_2093, n_2090, n_2091);
  nand g5276 (n_2062, n_2058, n_2059);
  or g5277 (n_1821, anoymous_7_126_n_47, b2);
  or g5278 (n_2438, n_1857, wc65);
  not gc65 (wc65, anoymous_7_126_n_47);
  nand g5280 (n_2059, anoymous_7_126_n_26, anoymous_7_126_n_47);
  or g5281 (n_1874, anoymous_7_126_n_47, b1);
  nand g5282 (n_1865, anoymous_7_126_n_47, b2);
  nand g5283 (n_2090, anoymous_7_126_n_47, n_1946);
  nand g5284 (anoymous_7_126_n_47, n_1964, a6);
  nand g5287 (n_1469, n_2040, n_2041);
  or g5288 (n_2041, anoymous_7_126_n_27, n_2039);
  or g5289 (n_2039, n_2037, wc66);
  not gc66 (wc66, a7);
  or g5291 (n_2037, wc67, anoymous_7_126_n_316);
  not gc67 (wc67, n_1856);
  or g5292 (anoymous_7_126_n_316, anoymous_7_126_n_29, n_2026);
  or g5293 (n_2026, n_1927, anoymous_7_126_n_28);
  nand g5294 (anoymous_7_126_n_322, anoymous_7_126_n_166, anoymous_7_126_n_202);
  or g5299 (n_2629, wc68, anoymous_7_126_n_200);
  not gc68 (wc68, n_1855);
  or g5300 (n_2630, n_1855, wc69);
  not gc69 (wc69, anoymous_7_126_n_200);
  nand g5301 (anoymous_7_126_n_30, n_2629, n_2630);
  nand g5302 (n_2425, n_2423, n_2424);
  nand g5303 (n_2063, n_2060, n_2061);
  nand g5304 (n_1946, n_1897, n_2023);
  nand g5306 (anoymous_7_126_n_200, n_1861, n_2020);
  nand g5307 (n_2631, n_1922, anoymous_7_126_n_181);
  or g5308 (n_2632, n_1922, anoymous_7_126_n_181);
  nand g5309 (anoymous_7_126_n_29, n_2631, n_2632);
  nand g5310 (n_2060, anoymous_7_126_n_27, anoymous_7_126_n_48);
  nand g5311 (n_2020, anoymous_7_126_n_162, anoymous_7_126_n_181);
  nand g5312 (n_2091, anoymous_7_126_n_48, b2);
  or g5313 (n_1921, anoymous_7_126_n_48, b2);
  nand g5314 (n_2023, anoymous_7_126_n_48, b1);
  nand g5319 (anoymous_7_126_n_48, n_2589, a7);
  or g5320 (n_2589, wc70, n_2587);
  not gc70 (wc70, n_2003);
  nand g5321 (n_2634, n_1919, anoymous_7_126_n_196);
  or g5322 (n_2635, n_1919, anoymous_7_126_n_196);
  nand g5323 (anoymous_7_126_n_28, n_2634, n_2635);
  or g5324 (anoymous_7_126_n_40, n_2011, b2);
  or g5325 (n_46, n_2017, b1);
  nand g5326 (n_2413, n_1858, n_2412);
  or g5327 (n_2011, n_2010, anoymous_7_126_n_152);
  nand g5328 (anoymous_7_126_n_643, n_1993, n_2416);
  nand g5330 (anoymous_7_126_n_511, n_1992, n_1993);
  nand g5331 (n_2286, n_2283, n_2284);
  or g5332 (n_2017, n_2016, b0);
  nand g5333 (anoymous_7_126_n_196, n_1857, n_1987);
  nand g5335 (n_2476, anoymous_7_126_n_25, n_1864);
  or g5336 (n_2636, wc71, n_1868);
  not gc71 (wc71, anoymous_7_126_n_340);
  or g5339 (n_2016, anoymous_7_126_n_156, n_1845);
  nand g5340 (n_2638, anoymous_7_126_n_340, anoymous_7_126_n_368);
  or g5341 (n_2639, anoymous_7_126_n_340, anoymous_7_126_n_368);
  nand g5342 (n_1967, n_2638, n_2639);
  nand g5343 (n_2640, n_1920, anoymous_7_126_n_167);
  or g5344 (n_2641, n_1920, anoymous_7_126_n_167);
  nand g5345 (anoymous_7_126_n_27, n_2640, n_2641);
  or g5346 (n_1992, wc72, b1);
  not gc72 (wc72, n_1876);
  nand g5347 (n_2283, n_1864, b1);
  or g5348 (n_2642, wc73, anoymous_7_126_n_193);
  not gc73 (wc73, n_1870);
  or g5349 (n_2643, n_1870, wc74);
  not gc74 (wc74, anoymous_7_126_n_193);
  nand g5350 (anoymous_7_126_n_26, n_2642, n_2643);
  or g5352 (n_2058, anoymous_7_126_n_340, wc75);
  not gc75 (wc75, n_1868);
  nand g5353 (anoymous_7_126_n_350, n_1975, n_2407);
  nand g5354 (n_1987, anoymous_7_126_n_156, anoymous_7_126_n_167);
  or g5355 (n_2010, n_1885, n_1835);
  nand g5356 (n_2644, anoymous_7_126_n_495, anoymous_7_126_n_672);
  or g5357 (n_2645, anoymous_7_126_n_495, anoymous_7_126_n_672);
  nand g5358 (n_1952, n_2644, n_2645);
  or g5359 (n_2284, n_1848, a0);
  nand g5360 (n_1951, anoymous_7_126_n_559, n_1981);
  or g5361 (n_2646, wc76, a3);
  not gc76 (wc76, anoymous_7_126_n_25);
  or g5362 (n_2647, anoymous_7_126_n_25, wc77);
  not gc77 (wc77, a3);
  nand g5363 (anoymous_7_126_n_672, n_2646, n_2647);
  or g5364 (n_2295, wc78, b1);
  not gc78 (wc78, n_1848);
  nand g5365 (n_1919, anoymous_7_126_n_152, n_1858);
  or g5366 (n_1931, n_1848, wc79);
  not gc79 (wc79, b1);
  nand g5367 (n_2648, anoymous_7_126_n_495, anoymous_7_126_n_536);
  or g5368 (n_2649, anoymous_7_126_n_495, anoymous_7_126_n_536);
  nand g5369 (n_1950, n_2648, n_2649);
  or g5370 (n_1845, anoymous_7_126_n_162, anoymous_7_126_n_166);
  nand g5371 (n_1864, n_1972, a1);
  nand g5372 (n_1922, anoymous_7_126_n_162, n_1861);
  nand g5373 (n_1993, anoymous_7_126_n_495, a3);
  nand g5374 (n_1920, anoymous_7_126_n_156, n_1857);
  nand g5375 (anoymous_7_126_n_368, n_1892, n_1975);
  or g5376 (n_2002, wc80, n_1856);
  not gc80 (wc80, n_1885);
  nand g5377 (n_1968, anoymous_7_126_n_388, n_1984);
  or g5378 (n_2061, wc81, a5);
  not gc81 (wc81, anoymous_7_126_n_25);
  nand g5379 (anoymous_7_126_n_193, n_1897, n_1978);
  nand g5380 (n_2407, anoymous_7_126_n_340, n_1892);
  nand g5381 (anoymous_7_126_n_167, n_1870, n_1897);
  or g5382 (n_2003, a7, wc82);
  not gc82 (wc82, b1);
  or g5383 (anoymous_7_126_n_559, a3, wc83);
  not gc83 (wc83, b0);
  or g5384 (anoymous_7_126_n_388, a5, wc84);
  not gc84 (wc84, b0);
  or g5385 (n_1972, a0, wc85);
  not gc85 (wc85, b0);
  or g5386 (anoymous_7_126_n_166, b6, b7);
  or g5387 (n_2650, wc86, b1);
  not gc86 (wc86, a3);
  or g5388 (n_2651, a3, wc87);
  not gc87 (wc87, b1);
  nand g5389 (anoymous_7_126_n_536, n_2650, n_2651);
  or g5390 (n_1981, wc88, b0);
  not gc88 (wc88, a3);
  nand g5391 (n_2424, b6, b5);
  or g5392 (n_1848, a1, wc89);
  not gc89 (wc89, b0);
  nand g5395 (anoymous_7_126_n_25, n_2652, n_2653);
  or g5396 (n_1984, wc90, b0);
  not gc90 (wc90, a5);
  or g5397 (n_1978, b2, b1);
  or g5398 (n_1975, wc91, b1);
  not gc91 (wc91, a5);
  nand g5399 (n_1897, b1, b2);
  or g5400 (anoymous_7_126_n_156, b2, b3);
  or g5401 (anoymous_7_126_n_152, b3, b4);
  or g5402 (anoymous_7_126_n_162, b4, b5);
  and g5403 (o7, n_46, wc92);
  not gc92 (wc92, anoymous_7_126_n_40);
  and g5404 (o6, n_46, n_1469);
  and g5406 (o4, n_1863, n_46);
  and g5408 (o2, n_1862, n_46);
  and g5409 (o1, wc93, n_46);
  not gc93 (wc93, anoymous_7_126_n_127);
  and g5410 (o0, n_1930, n_46);
  or g5412 (n_2652, wc94, b1);
  not gc94 (wc94, b0);
  or g5413 (n_2653, b0, wc95);
  not gc95 (wc95, b1);
  or g5415 (n_2416, anoymous_7_126_n_25, wc96);
  not gc96 (wc96, n_1876);
  or g5416 (n_2587, wc97, n_2016);
  not gc97 (wc97, n_2002);
  or g5417 (n_2412, wc98, n_1987);
  not gc98 (wc98, anoymous_7_126_n_152);
  or g5419 (n_2040, wc99, n_2589);
  not gc99 (wc99, anoymous_7_126_n_40);
  or g5420 (anoymous_7_126_n_181, n_2413, wc100);
  not gc100 (wc100, n_1857);
  or g5421 (n_2423, n_2020, wc101);
  not gc101 (wc101, n_1855);
  or g5422 (anoymous_7_126_n_202, n_2425, wc102);
  not gc102 (wc102, n_1861);
  or g5424 (anoymous_7_126_n_31, anoymous_7_126_n_166, anoymous_7_126_n_202);
  or g5426 (n_2625, wc103, n_1874);
  not gc103 (wc103, anoymous_7_126_n_388);
  or g5428 (n_2108, anoymous_7_126_n_64, n_2636);
  or g5429 (n_2440, wc104, n_2439);
  not gc104 (wc104, n_2438);
  or g5430 (n_1879, wc105, anoymous_7_126_n_61);
  not gc105 (wc105, anoymous_7_126_n_64);
  and g5431 (o5, n_46, wc106);
  not gc106 (wc106, anoymous_7_126_n_61);
  or g5432 (n_2122, n_2625, n_1879);
  or g5433 (n_2124, anoymous_7_126_n_47, wc107);
  not gc107 (wc107, anoymous_7_126_n_59);
  or g5434 (anoymous_7_126_n_62, wc108, anoymous_7_126_n_59);
  not gc108 (wc108, anoymous_7_126_n_61);
  or g5435 (anoymous_7_126_n_71, anoymous_7_126_n_48, wc109);
  not gc109 (wc109, anoymous_7_126_n_59);
  or g5436 (anoymous_7_126_n_70, wc110, n_2125);
  not gc110 (wc110, n_2124);
  or g5437 (n_1889, anoymous_7_126_n_27, wc111);
  not gc111 (wc111, anoymous_7_126_n_69);
  or g5438 (n_2131, wc112, anoymous_7_126_n_69);
  not gc112 (wc112, anoymous_7_126_n_27);
  or g5439 (n_2146, anoymous_7_126_n_26, wc113);
  not gc113 (wc113, anoymous_7_126_n_68);
  or g5440 (n_1893, wc114, anoymous_7_126_n_68);
  not gc114 (wc114, anoymous_7_126_n_26);
  or g5442 (n_2448, wc115, anoymous_7_126_n_675);
  not gc115 (wc115, n_1889);
  or g5443 (anoymous_7_126_n_658, wc116, n_2449);
  not gc116 (wc116, n_2131);
  or g5444 (n_2604, wc117, n_1820);
  not gc117 (wc117, anoymous_7_126_n_589);
  or g5445 (n_2171, wc118, n_2169);
  not gc118 (wc118, anoymous_7_126_n_658);
  or g5447 (n_2246, wc119, anoymous_7_126_n_93);
  not gc119 (wc119, n_1961);
  or g5448 (n_2197, wc120, n_2196);
  not gc120 (wc120, n_2195);
  or g5449 (n_2228, wc121, anoymous_7_126_n_93);
  not gc121 (wc121, n_1952);
  or g5450 (n_2210, wc122, anoymous_7_126_n_93);
  not gc122 (wc122, n_1955);
  or g5451 (anoymous_7_126_n_102, anoymous_7_126_n_71, wc123);
  not gc123 (wc123, anoymous_7_126_n_89);
  or g5452 (anoymous_7_126_n_94, wc124, anoymous_7_126_n_90);
  not gc124 (wc124, anoymous_7_126_n_93);
  or g5453 (anoymous_7_126_n_91, anoymous_7_126_n_89, wc125);
  not gc125 (wc125, anoymous_7_126_n_90);
  and g5454 (o3, n_46, wc126);
  not gc126 (wc126, anoymous_7_126_n_90);
  or g5455 (n_2260, n_2604, anoymous_7_126_n_94);
  or g5456 (n_1849, wc127, anoymous_7_126_n_100);
  not gc127 (wc127, anoymous_7_126_n_29);
  or g5457 (n_1871, wc128, anoymous_7_126_n_98);
  not gc128 (wc128, anoymous_7_126_n_27);
  or g5458 (n_1929, wc129, anoymous_7_126_n_101);
  not gc129 (wc129, anoymous_7_126_n_30);
  or g5459 (n_2381, anoymous_7_126_n_166, wc130);
  not gc130 (wc130, anoymous_7_126_n_101);
  or g5460 (n_1852, anoymous_7_126_n_102, wc131);
  not gc131 (wc131, anoymous_7_126_n_101);
  or g5461 (n_1905, wc132, anoymous_7_126_n_101);
  not gc132 (wc132, anoymous_7_126_n_102);
  or g5462 (n_2353, anoymous_7_126_n_27, wc133);
  not gc133 (wc133, anoymous_7_126_n_98);
  or g5463 (n_2398, anoymous_7_126_n_29, wc134);
  not gc134 (wc134, anoymous_7_126_n_100);
  or g5464 (n_2477, wc135, anoymous_7_126_n_97);
  not gc135 (wc135, anoymous_7_126_n_26);
  or g5465 (anoymous_7_126_n_723, n_2287, wc136);
  not gc136 (wc136, n_1873);
  or g5466 (n_2320, wc137, n_1917);
  not gc137 (wc137, anoymous_7_126_n_99);
  or g5467 (n_2479, wc138, n_2478);
  not gc138 (wc138, n_2284);
  or g5468 (anoymous_7_126_n_879, n_2479, wc139);
  not gc139 (wc139, n_1871);
  or g5469 (anoymous_7_126_n_734, wc140, n_2335);
  not gc140 (wc140, n_2334);
  or g5470 (anoymous_7_126_n_821, wc141, anoymous_7_126_n_809);
  not gc141 (wc141, n_1935);
  or g5471 (n_2384, anoymous_7_126_n_732, wc142);
  not gc142 (wc142, n_2380);
  or g5472 (n_2386, n_2384, wc143);
  not gc143 (wc143, n_2383);
  or g5473 (anoymous_7_126_n_127, b7, wc144);
  not gc144 (wc144, n_2401);
endmodule

