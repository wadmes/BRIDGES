
module test ( a_0, a_1, a_2, a_3, b_0, b_1, b_2, b_3, sum_0, sum_1, sum_2, sum_3, sum_4, sum_5, sum_6, sum_7);
  input a_0;
  input a_1;
  input a_2;
  input a_3;

  input b_0;
  input b_1;
  input b_2;
  input b_3;

  output sum_0;
  output sum_1;
  output sum_2;
  output sum_3;
  output sum_4;
  output sum_5;
  output sum_6;
  output sum_7;

	not gate_mult_9_n65 (mult_9_n65, a_0);
	not gate_mult_9_n64 (mult_9_n64, a_1);
	not gate_mult_9_n63 (mult_9_n63, a_2);
	not gate_mult_9_n62 (mult_9_n62, a_3);
	not gate_mult_9_n61 (mult_9_n61, b_0);
	not gate_mult_9_n60 (mult_9_n60, b_1);
	not gate_mult_9_n59 (mult_9_n59, b_2);
	not gate_mult_9_n58 (mult_9_n58, b_3);
	nor gate_sum_0 (sum_0, mult_9_n65, mult_9_n61);
	nor gate_mult_9_n57 (mult_9_n57, mult_9_n65, mult_9_n60);
	nor gate_mult_9_n56 (mult_9_n56, mult_9_n65, mult_9_n59);
	nor gate_mult_9_n55 (mult_9_n55, mult_9_n65, mult_9_n58);
	nor gate_mult_9_n54 (mult_9_n54, mult_9_n64, mult_9_n61);
	nor gate_mult_9_n53 (mult_9_n53, mult_9_n64, mult_9_n60);
	nor gate_mult_9_n52 (mult_9_n52, mult_9_n64, mult_9_n59);
	nor gate_mult_9_n51 (mult_9_n51, mult_9_n64, mult_9_n58);
	nor gate_mult_9_n50 (mult_9_n50, mult_9_n63, mult_9_n61);
	nor gate_mult_9_n49 (mult_9_n49, mult_9_n63, mult_9_n60);
	nor gate_mult_9_n48 (mult_9_n48, mult_9_n63, mult_9_n59);
	nor gate_mult_9_n47 (mult_9_n47, mult_9_n63, mult_9_n58);
	nor gate_mult_9_n46 (mult_9_n46, mult_9_n62, mult_9_n61);
	nor gate_mult_9_n45 (mult_9_n45, mult_9_n62, mult_9_n60);
	nor gate_mult_9_n44 (mult_9_n44, mult_9_n62, mult_9_n59);
	nor gate_mult_9_n43 (mult_9_n43, mult_9_n62, mult_9_n58);
	and gate_mult_9_n41 (mult_9_n41, mult_9_n53, mult_9_n56);
	xor gate_mult_9_n42 (mult_9_n42, mult_9_n56, mult_9_n53);
	and gate_mult_9_n39 (mult_9_n39, mult_9_n46, mult_9_n49);
	xor gate_mult_9_n40 (mult_9_n40, mult_9_n49, mult_9_n46);
	xor gate_mult_9_n36 (mult_9_n36, mult_9_n55, mult_9_n52);
	and gate_mult_9_n35 (mult_9_n35, mult_9_n52, mult_9_n55);
	and gate_mult_9_n34 (mult_9_n34, mult_9_n36, mult_9_n41);
	or gate_mult_9_n37 (mult_9_n37, mult_9_n35, mult_9_n34);
	xor gate_mult_9_n38 (mult_9_n38, mult_9_n41, mult_9_n36);
	and gate_mult_9_n32 (mult_9_n32, mult_9_n45, mult_9_n51);
	xor gate_mult_9_n33 (mult_9_n33, mult_9_n51, mult_9_n45);
	xor gate_mult_9_n29 (mult_9_n29, mult_9_n48, mult_9_n39);
	and gate_mult_9_n28 (mult_9_n28, mult_9_n39, mult_9_n48);
	and gate_mult_9_n27 (mult_9_n27, mult_9_n29, mult_9_n33);
	or gate_mult_9_n30 (mult_9_n30, mult_9_n28, mult_9_n27);
	xor gate_mult_9_n31 (mult_9_n31, mult_9_n33, mult_9_n29);
	xor gate_mult_9_n24 (mult_9_n24, mult_9_n47, mult_9_n44);
	and gate_mult_9_n23 (mult_9_n23, mult_9_n44, mult_9_n47);
	and gate_mult_9_n22 (mult_9_n22, mult_9_n24, mult_9_n32);
	or gate_mult_9_n25 (mult_9_n25, mult_9_n23, mult_9_n22);
	xor gate_mult_9_n26 (mult_9_n26, mult_9_n32, mult_9_n24);
	and gate_mult_9_n21 (mult_9_n21, mult_9_n57, mult_9_n54);
	xor gate_sum_1 (sum_1, mult_9_n54, mult_9_n57);
	xor gate_mult_9_n15 (mult_9_n15, mult_9_n50, mult_9_n42);
	and gate_mult_9_n14 (mult_9_n14, mult_9_n42, mult_9_n50);
	and gate_mult_9_n13 (mult_9_n13, mult_9_n15, mult_9_n21);
	or gate_mult_9_n20 (mult_9_n20, mult_9_n14, mult_9_n13);
	xor gate_sum_2 (sum_2, mult_9_n21, mult_9_n15);
	xor gate_mult_9_n12 (mult_9_n12, mult_9_n40, mult_9_n38);
	and gate_mult_9_n11 (mult_9_n11, mult_9_n38, mult_9_n40);
	and gate_mult_9_n10 (mult_9_n10, mult_9_n12, mult_9_n20);
	or gate_mult_9_n19 (mult_9_n19, mult_9_n11, mult_9_n10);
	xor gate_sum_3 (sum_3, mult_9_n20, mult_9_n12);
	xor gate_mult_9_n9 (mult_9_n9, mult_9_n37, mult_9_n31);
	and gate_mult_9_n8 (mult_9_n8, mult_9_n31, mult_9_n37);
	and gate_mult_9_n7 (mult_9_n7, mult_9_n19, mult_9_n9);
	or gate_mult_9_n18 (mult_9_n18, mult_9_n8, mult_9_n7);
	xor gate_sum_4 (sum_4, mult_9_n9, mult_9_n19);
	xor gate_mult_9_n6 (mult_9_n6, mult_9_n26, mult_9_n30);
	and gate_mult_9_n5 (mult_9_n5, mult_9_n30, mult_9_n26);
	and gate_mult_9_n4 (mult_9_n4, mult_9_n18, mult_9_n6);
	or gate_mult_9_n17 (mult_9_n17, mult_9_n5, mult_9_n4);
	xor gate_sum_5 (sum_5, mult_9_n6, mult_9_n18);
	xor gate_mult_9_n3 (mult_9_n3, mult_9_n43, mult_9_n25);
	and gate_mult_9_n2 (mult_9_n2, mult_9_n25, mult_9_n43);
	and gate_mult_9_n1 (mult_9_n1, mult_9_n17, mult_9_n3);
	or gate_mult_9_n16 (mult_9_n16, mult_9_n2, mult_9_n1);
	xor gate_sum_6 (sum_6, mult_9_n3, mult_9_n17);
	buf gate_sum_7 (sum_7, mult_9_n16);
endmodule

