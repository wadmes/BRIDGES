module test (a3, a2, a1, a0, b3, b2, b1, b0, o3, o2, o1, o0);
  input a3, a2, a1, a0, b3, b2, b1, b0;
  output o3, o2, o1, o0;
  wire a3, a2, a1, a0, b3, b2, b1, b0;
  wire o3, o2, o1, o0;
  wire n_244, n_247, n_250, n_266, n_268, n_275, n_279, n_286;
  wire n_288, n_289, n_292, n_303, n_319, n_320, n_322, n_330;
  wire n_331, n_336, n_338, n_339, n_340, n_341, n_342, n_343;
  wire n_344, n_345, n_346, n_347, n_348, n_355, n_356, n_357;
  wire n_360, n_363, n_366, n_373, n_374, n_375, n_378, n_385;
  wire n_386, n_387, n_390, n_393, n_396, n_399, n_406, n_407;
  wire n_408, n_413, n_414, n_417, n_420, n_427, n_428, n_429;
  wire n_446, n_447, n_448, n_449, n_450, n_451, n_452, n_453;
  wire n_462, n_463, n_464, n_465, n_468, n_489, n_490, n_491;
  wire n_492, n_493, n_494, n_495, n_496, n_497, n_498, n_507;
  wire n_508, n_509, n_510;
  or g306 (n_250, b1, wc);
  not gc (wc, a2);
  or g478 (n_320, wc0, a1);
  not gc0 (wc0, b0);
  nand g569 (n_341, n_250, b2);
  or g583 (n_348, a3, wc1);
  not gc1 (wc1, b3);
  or g699 (o0, n_497, n_498);
  or g700 (n_498, n_495, n_496);
  nand g701 (n_495, n_286, n_292);
  or g702 (n_497, wc2, n_494);
  not gc2 (wc2, n_493);
  nand g703 (n_494, n_289, n_275);
  or g704 (o1, n_452, n_453);
  nand g705 (n_496, n_491, n_492);
  or g706 (n_286, n_468, a3);
  nand g707 (n_453, n_450, n_451);
  or g708 (n_275, n_420, wc3);
  not gc3 (wc3, a1);
  or g709 (n_468, wc4, b3);
  not gc4 (wc4, n_344);
  or g710 (n_492, wc5, n_322);
  not gc5 (wc5, n_347);
  or g711 (n_347, wc6, n_465);
  not gc6 (wc6, n_464);
  nand g712 (n_420, n_342, a0);
  or g713 (n_451, n_447, wc7);
  not gc7 (wc7, a2);
  nand g714 (n_344, n_428, n_429);
  nand g715 (n_491, n_348, n_268);
  nand g716 (n_447, n_336, a1);
  or g717 (n_450, n_446, a2);
  nand g718 (n_452, n_448, n_449);
  nand g719 (n_342, n_407, n_408);
  nand g720 (n_268, n_386, n_387);
  or g721 (o2, wc8, n_510);
  not gc8 (wc8, n_509);
  nand g722 (n_428, n_343, a2);
  nand g723 (n_465, n_462, n_463);
  or g724 (n_292, n_417, a2);
  or g725 (n_463, wc9, b2);
  not gc9 (wc9, n_338);
  or g726 (n_408, n_406, wc10);
  not gc10 (wc10, b0);
  nand g727 (n_336, n_393, n_288);
  or g728 (n_289, n_390, wc11);
  not gc11 (wc11, n_250);
  or g729 (n_493, n_490, a2);
  nand g730 (n_510, n_507, n_508);
  or g731 (n_446, n_247, wc12);
  not gc12 (wc12, b1);
  nand g732 (n_449, n_345, n_303);
  or g733 (n_343, n_266, wc13);
  not gc13 (wc13, n_414);
  or g734 (n_509, n_247, wc14);
  not gc14 (wc14, a2);
  or g735 (n_429, n_427, wc15);
  not gc15 (wc15, b2);
  nand g736 (n_417, n_340, b1);
  or g737 (n_386, wc16, b2);
  not gc16 (wc16, n_266);
  nand g740 (n_462, n_339, a1);
  or g741 (n_387, n_385, b0);
  nand g742 (n_427, n_279, a1);
  or g743 (n_414, n_413, wc17);
  not gc17 (wc17, b1);
  nand g744 (n_303, n_356, n_357);
  or g745 (n_448, wc18, n_288);
  not gc18 (wc18, n_346);
  or g746 (n_508, n_250, n_319);
  nand g747 (n_406, n_341, a3);
  or g748 (n_407, n_319, a2);
  nand g749 (n_340, n_288, n_399);
  nand g750 (n_266, n_374, n_375);
  or g751 (n_339, wc19, n_279);
  not gc19 (wc19, n_396);
  or g752 (n_338, wc20, a2);
  not gc20 (wc20, n_360);
  or g753 (n_247, n_378, wc21);
  not gc21 (wc21, b0);
  or g754 (n_393, n_319, a3);
  or g755 (n_507, n_378, n_330);
  or g756 (n_390, n_288, n_320);
  or g757 (n_490, n_489, wc22);
  not gc22 (wc22, a0);
  nand g758 (n_345, n_244, n_331);
  or g759 (n_413, n_320, b2);
  or g760 (n_288, wc23, n_244);
  not gc23 (wc23, b2);
  or g761 (n_399, n_244, wc24);
  not gc24 (wc24, a1);
  or g762 (n_378, n_244, b2);
  or g763 (n_464, n_250, wc25);
  not gc25 (wc25, a0);
  or g764 (n_489, n_320, n_244);
  or g765 (n_385, n_250, wc26);
  not gc26 (wc26, b2);
  or g766 (n_375, n_373, wc27);
  not gc27 (wc27, b0);
  or g767 (n_374, n_330, wc28);
  not gc28 (wc28, a1);
  nand g768 (n_279, n_250, n_366);
  or g769 (n_356, n_330, wc29);
  not gc29 (wc29, a2);
  nand g770 (n_346, n_250, n_363);
  or g771 (n_319, n_331, wc30);
  not gc30 (wc30, b0);
  or g772 (n_360, wc31, b1);
  not gc31 (wc31, n_320);
  or g773 (n_357, n_355, wc32);
  not gc32 (wc32, b0);
  or g774 (n_355, wc33, b1);
  not gc33 (wc33, a1);
  or g775 (n_331, b3, b2);
  or g776 (n_330, wc34, b0);
  not gc34 (wc34, b1);
  nand g777 (n_322, b3, a3);
  or g778 (n_363, b1, b0);
  nand g779 (n_366, a2, a0);
  or g780 (n_373, wc35, b1);
  not gc35 (wc35, a0);
  or g781 (n_396, wc36, b0);
  not gc36 (wc36, a2);
  or g782 (n_244, wc37, b3);
  not gc37 (wc37, a3);
  nor g783 (o3, n_247, b1);
endmodule

