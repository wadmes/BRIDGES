
module test ( a_0, a_1, a_2, a_3, a_4, a_5, a_6, a_7, b_0, b_1, b_2, b_3, b_4, b_5, b_6, b_7, 
  sum_0, sum_1, sum_2, sum_3, sum_4, sum_5, sum_6, sum_7, sum_8, sum_9, sum_10, sum_11, 
   sum_12, sum_13, sum_14, sum_15);
  
  input a_0;
  input a_1;
  input a_2;
  input a_3;
  input a_4;
  input a_5;
  input a_6;
  input a_7;

  input b_0;
  input b_1;
  input b_2;
  input b_3;
  input b_4;
  input b_5;
  input b_6;
  input b_7;
  
  output sum_0;
  output sum_1;
  output sum_2;
  output sum_3;
  output sum_4;
  output sum_5;
  output sum_6;
  output sum_7;
  output sum_8;
  output sum_9;
  output sum_10;
  output sum_11;
  output sum_12;
  output sum_13;
  output sum_14;
  output sum_15;
 

	not gate_mult_9_n321 (mult_9_n321, a_0);
	not gate_mult_9_n320 (mult_9_n320, a_1);
	not gate_mult_9_n319 (mult_9_n319, a_2);
	not gate_mult_9_n318 (mult_9_n318, a_3);
	not gate_mult_9_n317 (mult_9_n317, a_4);
	not gate_mult_9_n316 (mult_9_n316, a_5);
	not gate_mult_9_n315 (mult_9_n315, a_6);
	not gate_mult_9_n314 (mult_9_n314, a_7);
	not gate_mult_9_n313 (mult_9_n313, b_0);
	not gate_mult_9_n312 (mult_9_n312, b_1);
	not gate_mult_9_n311 (mult_9_n311, b_2);
	not gate_mult_9_n310 (mult_9_n310, b_3);
	not gate_mult_9_n309 (mult_9_n309, b_4);
	not gate_mult_9_n308 (mult_9_n308, b_5);
	not gate_mult_9_n307 (mult_9_n307, b_6);
	not gate_mult_9_n306 (mult_9_n306, b_7);
	nor gate_sum_0 (sum_0, mult_9_n321, mult_9_n313);
	nor gate_mult_9_n305 (mult_9_n305, mult_9_n321, mult_9_n312);
	nor gate_mult_9_n304 (mult_9_n304, mult_9_n321, mult_9_n311);
	nor gate_mult_9_n303 (mult_9_n303, mult_9_n321, mult_9_n310);
	nor gate_mult_9_n302 (mult_9_n302, mult_9_n321, mult_9_n309);
	nor gate_mult_9_n301 (mult_9_n301, mult_9_n321, mult_9_n308);
	nor gate_mult_9_n300 (mult_9_n300, mult_9_n321, mult_9_n307);
	nor gate_mult_9_n299 (mult_9_n299, mult_9_n321, mult_9_n306);
	nor gate_mult_9_n298 (mult_9_n298, mult_9_n320, mult_9_n313);
	nor gate_mult_9_n297 (mult_9_n297, mult_9_n320, mult_9_n312);
	nor gate_mult_9_n296 (mult_9_n296, mult_9_n320, mult_9_n311);
	nor gate_mult_9_n295 (mult_9_n295, mult_9_n320, mult_9_n310);
	nor gate_mult_9_n294 (mult_9_n294, mult_9_n320, mult_9_n309);
	nor gate_mult_9_n293 (mult_9_n293, mult_9_n320, mult_9_n308);
	nor gate_mult_9_n292 (mult_9_n292, mult_9_n320, mult_9_n307);
	nor gate_mult_9_n291 (mult_9_n291, mult_9_n320, mult_9_n306);
	nor gate_mult_9_n290 (mult_9_n290, mult_9_n319, mult_9_n313);
	nor gate_mult_9_n289 (mult_9_n289, mult_9_n319, mult_9_n312);
	nor gate_mult_9_n288 (mult_9_n288, mult_9_n319, mult_9_n311);
	nor gate_mult_9_n287 (mult_9_n287, mult_9_n319, mult_9_n310);
	nor gate_mult_9_n286 (mult_9_n286, mult_9_n319, mult_9_n309);
	nor gate_mult_9_n285 (mult_9_n285, mult_9_n319, mult_9_n308);
	nor gate_mult_9_n284 (mult_9_n284, mult_9_n319, mult_9_n307);
	nor gate_mult_9_n283 (mult_9_n283, mult_9_n319, mult_9_n306);
	nor gate_mult_9_n282 (mult_9_n282, mult_9_n318, mult_9_n313);
	nor gate_mult_9_n281 (mult_9_n281, mult_9_n318, mult_9_n312);
	nor gate_mult_9_n280 (mult_9_n280, mult_9_n318, mult_9_n311);
	nor gate_mult_9_n279 (mult_9_n279, mult_9_n318, mult_9_n310);
	nor gate_mult_9_n278 (mult_9_n278, mult_9_n318, mult_9_n309);
	nor gate_mult_9_n277 (mult_9_n277, mult_9_n318, mult_9_n308);
	nor gate_mult_9_n276 (mult_9_n276, mult_9_n318, mult_9_n307);
	nor gate_mult_9_n275 (mult_9_n275, mult_9_n318, mult_9_n306);
	nor gate_mult_9_n274 (mult_9_n274, mult_9_n317, mult_9_n313);
	nor gate_mult_9_n273 (mult_9_n273, mult_9_n317, mult_9_n312);
	nor gate_mult_9_n272 (mult_9_n272, mult_9_n317, mult_9_n311);
	nor gate_mult_9_n271 (mult_9_n271, mult_9_n317, mult_9_n310);
	nor gate_mult_9_n270 (mult_9_n270, mult_9_n317, mult_9_n309);
	nor gate_mult_9_n269 (mult_9_n269, mult_9_n317, mult_9_n308);
	nor gate_mult_9_n268 (mult_9_n268, mult_9_n317, mult_9_n307);
	nor gate_mult_9_n267 (mult_9_n267, mult_9_n317, mult_9_n306);
	nor gate_mult_9_n266 (mult_9_n266, mult_9_n316, mult_9_n313);
	nor gate_mult_9_n265 (mult_9_n265, mult_9_n316, mult_9_n312);
	nor gate_mult_9_n264 (mult_9_n264, mult_9_n316, mult_9_n311);
	nor gate_mult_9_n263 (mult_9_n263, mult_9_n316, mult_9_n310);
	nor gate_mult_9_n262 (mult_9_n262, mult_9_n316, mult_9_n309);
	nor gate_mult_9_n261 (mult_9_n261, mult_9_n316, mult_9_n308);
	nor gate_mult_9_n260 (mult_9_n260, mult_9_n316, mult_9_n307);
	nor gate_mult_9_n259 (mult_9_n259, mult_9_n316, mult_9_n306);
	nor gate_mult_9_n258 (mult_9_n258, mult_9_n315, mult_9_n313);
	nor gate_mult_9_n257 (mult_9_n257, mult_9_n315, mult_9_n312);
	nor gate_mult_9_n256 (mult_9_n256, mult_9_n315, mult_9_n311);
	nor gate_mult_9_n255 (mult_9_n255, mult_9_n315, mult_9_n310);
	nor gate_mult_9_n254 (mult_9_n254, mult_9_n315, mult_9_n309);
	nor gate_mult_9_n253 (mult_9_n253, mult_9_n315, mult_9_n308);
	nor gate_mult_9_n252 (mult_9_n252, mult_9_n315, mult_9_n307);
	nor gate_mult_9_n251 (mult_9_n251, mult_9_n315, mult_9_n306);
	nor gate_mult_9_n250 (mult_9_n250, mult_9_n314, mult_9_n313);
	nor gate_mult_9_n249 (mult_9_n249, mult_9_n314, mult_9_n312);
	nor gate_mult_9_n248 (mult_9_n248, mult_9_n314, mult_9_n311);
	nor gate_mult_9_n247 (mult_9_n247, mult_9_n314, mult_9_n310);
	nor gate_mult_9_n246 (mult_9_n246, mult_9_n314, mult_9_n309);
	nor gate_mult_9_n245 (mult_9_n245, mult_9_n314, mult_9_n308);
	nor gate_mult_9_n244 (mult_9_n244, mult_9_n314, mult_9_n307);
	nor gate_mult_9_n243 (mult_9_n243, mult_9_n314, mult_9_n306);
	and gate_mult_9_n241 (mult_9_n241, mult_9_n297, mult_9_n304);
	xor gate_mult_9_n242 (mult_9_n242, mult_9_n304, mult_9_n297);
	and gate_mult_9_n239 (mult_9_n239, mult_9_n282, mult_9_n289);
	xor gate_mult_9_n240 (mult_9_n240, mult_9_n289, mult_9_n282);
	xor gate_mult_9_n236 (mult_9_n236, mult_9_n303, mult_9_n296);
	and gate_mult_9_n235 (mult_9_n235, mult_9_n296, mult_9_n303);
	and gate_mult_9_n234 (mult_9_n234, mult_9_n236, mult_9_n241);
	or gate_mult_9_n237 (mult_9_n237, mult_9_n235, mult_9_n234);
	xor gate_mult_9_n238 (mult_9_n238, mult_9_n241, mult_9_n236);
	and gate_mult_9_n232 (mult_9_n232, mult_9_n274, mult_9_n281);
	xor gate_mult_9_n233 (mult_9_n233, mult_9_n281, mult_9_n274);
	xor gate_mult_9_n229 (mult_9_n229, mult_9_n302, mult_9_n295);
	and gate_mult_9_n228 (mult_9_n228, mult_9_n295, mult_9_n302);
	and gate_mult_9_n227 (mult_9_n227, mult_9_n229, mult_9_n288);
	or gate_mult_9_n230 (mult_9_n230, mult_9_n228, mult_9_n227);
	xor gate_mult_9_n231 (mult_9_n231, mult_9_n288, mult_9_n229);
	xor gate_mult_9_n224 (mult_9_n224, mult_9_n239, mult_9_n233);
	and gate_mult_9_n223 (mult_9_n223, mult_9_n233, mult_9_n239);
	and gate_mult_9_n222 (mult_9_n222, mult_9_n224, mult_9_n237);
	or gate_mult_9_n225 (mult_9_n225, mult_9_n223, mult_9_n222);
	xor gate_mult_9_n226 (mult_9_n226, mult_9_n237, mult_9_n224);
	and gate_mult_9_n220 (mult_9_n220, mult_9_n266, mult_9_n273);
	xor gate_mult_9_n221 (mult_9_n221, mult_9_n273, mult_9_n266);
	xor gate_mult_9_n217 (mult_9_n217, mult_9_n301, mult_9_n294);
	and gate_mult_9_n216 (mult_9_n216, mult_9_n294, mult_9_n301);
	and gate_mult_9_n215 (mult_9_n215, mult_9_n217, mult_9_n287);
	or gate_mult_9_n218 (mult_9_n218, mult_9_n216, mult_9_n215);
	xor gate_mult_9_n219 (mult_9_n219, mult_9_n287, mult_9_n217);
	xor gate_mult_9_n212 (mult_9_n212, mult_9_n280, mult_9_n232);
	and gate_mult_9_n211 (mult_9_n211, mult_9_n232, mult_9_n280);
	and gate_mult_9_n210 (mult_9_n210, mult_9_n212, mult_9_n221);
	or gate_mult_9_n213 (mult_9_n213, mult_9_n211, mult_9_n210);
	xor gate_mult_9_n214 (mult_9_n214, mult_9_n221, mult_9_n212);
	xor gate_mult_9_n207 (mult_9_n207, mult_9_n230, mult_9_n219);
	and gate_mult_9_n206 (mult_9_n206, mult_9_n219, mult_9_n230);
	and gate_mult_9_n205 (mult_9_n205, mult_9_n207, mult_9_n214);
	or gate_mult_9_n208 (mult_9_n208, mult_9_n206, mult_9_n205);
	xor gate_mult_9_n209 (mult_9_n209, mult_9_n214, mult_9_n207);
	and gate_mult_9_n203 (mult_9_n203, mult_9_n258, mult_9_n265);
	xor gate_mult_9_n204 (mult_9_n204, mult_9_n265, mult_9_n258);
	xor gate_mult_9_n200 (mult_9_n200, mult_9_n300, mult_9_n293);
	and gate_mult_9_n199 (mult_9_n199, mult_9_n293, mult_9_n300);
	and gate_mult_9_n198 (mult_9_n198, mult_9_n200, mult_9_n272);
	or gate_mult_9_n201 (mult_9_n201, mult_9_n199, mult_9_n198);
	xor gate_mult_9_n202 (mult_9_n202, mult_9_n272, mult_9_n200);
	xor gate_mult_9_n195 (mult_9_n195, mult_9_n286, mult_9_n279);
	and gate_mult_9_n194 (mult_9_n194, mult_9_n279, mult_9_n286);
	and gate_mult_9_n193 (mult_9_n193, mult_9_n195, mult_9_n220);
	or gate_mult_9_n196 (mult_9_n196, mult_9_n194, mult_9_n193);
	xor gate_mult_9_n197 (mult_9_n197, mult_9_n220, mult_9_n195);
	xor gate_mult_9_n190 (mult_9_n190, mult_9_n204, mult_9_n218);
	and gate_mult_9_n189 (mult_9_n189, mult_9_n218, mult_9_n204);
	and gate_mult_9_n188 (mult_9_n188, mult_9_n190, mult_9_n197);
	or gate_mult_9_n191 (mult_9_n191, mult_9_n189, mult_9_n188);
	xor gate_mult_9_n192 (mult_9_n192, mult_9_n197, mult_9_n190);
	xor gate_mult_9_n185 (mult_9_n185, mult_9_n202, mult_9_n213);
	and gate_mult_9_n184 (mult_9_n184, mult_9_n213, mult_9_n202);
	and gate_mult_9_n183 (mult_9_n183, mult_9_n208, mult_9_n185);
	or gate_mult_9_n186 (mult_9_n186, mult_9_n184, mult_9_n183);
	xor gate_mult_9_n187 (mult_9_n187, mult_9_n185, mult_9_n208);
	and gate_mult_9_n181 (mult_9_n181, mult_9_n250, mult_9_n257);
	xor gate_mult_9_n182 (mult_9_n182, mult_9_n257, mult_9_n250);
	xor gate_mult_9_n178 (mult_9_n178, mult_9_n299, mult_9_n292);
	and gate_mult_9_n177 (mult_9_n177, mult_9_n292, mult_9_n299);
	and gate_mult_9_n176 (mult_9_n176, mult_9_n178, mult_9_n271);
	or gate_mult_9_n179 (mult_9_n179, mult_9_n177, mult_9_n176);
	xor gate_mult_9_n180 (mult_9_n180, mult_9_n271, mult_9_n178);
	xor gate_mult_9_n173 (mult_9_n173, mult_9_n264, mult_9_n278);
	and gate_mult_9_n172 (mult_9_n172, mult_9_n278, mult_9_n264);
	and gate_mult_9_n171 (mult_9_n171, mult_9_n173, mult_9_n285);
	or gate_mult_9_n174 (mult_9_n174, mult_9_n172, mult_9_n171);
	xor gate_mult_9_n175 (mult_9_n175, mult_9_n285, mult_9_n173);
	xor gate_mult_9_n168 (mult_9_n168, mult_9_n203, mult_9_n182);
	and gate_mult_9_n167 (mult_9_n167, mult_9_n182, mult_9_n203);
	and gate_mult_9_n166 (mult_9_n166, mult_9_n168, mult_9_n201);
	or gate_mult_9_n169 (mult_9_n169, mult_9_n167, mult_9_n166);
	xor gate_mult_9_n170 (mult_9_n170, mult_9_n201, mult_9_n168);
	xor gate_mult_9_n163 (mult_9_n163, mult_9_n196, mult_9_n175);
	and gate_mult_9_n162 (mult_9_n162, mult_9_n175, mult_9_n196);
	and gate_mult_9_n161 (mult_9_n161, mult_9_n163, mult_9_n180);
	or gate_mult_9_n164 (mult_9_n164, mult_9_n162, mult_9_n161);
	xor gate_mult_9_n165 (mult_9_n165, mult_9_n180, mult_9_n163);
	xor gate_mult_9_n158 (mult_9_n158, mult_9_n170, mult_9_n191);
	and gate_mult_9_n157 (mult_9_n157, mult_9_n191, mult_9_n170);
	and gate_mult_9_n156 (mult_9_n156, mult_9_n158, mult_9_n165);
	or gate_mult_9_n159 (mult_9_n159, mult_9_n157, mult_9_n156);
	xor gate_mult_9_n160 (mult_9_n160, mult_9_n165, mult_9_n158);
	and gate_mult_9_n154 (mult_9_n154, mult_9_n249, mult_9_n256);
	xor gate_mult_9_n155 (mult_9_n155, mult_9_n256, mult_9_n249);
	xor gate_mult_9_n151 (mult_9_n151, mult_9_n270, mult_9_n277);
	and gate_mult_9_n150 (mult_9_n150, mult_9_n277, mult_9_n270);
	and gate_mult_9_n149 (mult_9_n149, mult_9_n151, mult_9_n263);
	or gate_mult_9_n152 (mult_9_n152, mult_9_n150, mult_9_n149);
	xor gate_mult_9_n153 (mult_9_n153, mult_9_n263, mult_9_n151);
	xor gate_mult_9_n146 (mult_9_n146, mult_9_n291, mult_9_n284);
	and gate_mult_9_n145 (mult_9_n145, mult_9_n284, mult_9_n291);
	and gate_mult_9_n144 (mult_9_n144, mult_9_n146, mult_9_n181);
	or gate_mult_9_n147 (mult_9_n147, mult_9_n145, mult_9_n144);
	xor gate_mult_9_n148 (mult_9_n148, mult_9_n181, mult_9_n146);
	xor gate_mult_9_n141 (mult_9_n141, mult_9_n155, mult_9_n179);
	and gate_mult_9_n140 (mult_9_n140, mult_9_n179, mult_9_n155);
	and gate_mult_9_n139 (mult_9_n139, mult_9_n141, mult_9_n174);
	or gate_mult_9_n142 (mult_9_n142, mult_9_n140, mult_9_n139);
	xor gate_mult_9_n143 (mult_9_n143, mult_9_n174, mult_9_n141);
	xor gate_mult_9_n136 (mult_9_n136, mult_9_n148, mult_9_n153);
	and gate_mult_9_n135 (mult_9_n135, mult_9_n153, mult_9_n148);
	and gate_mult_9_n134 (mult_9_n134, mult_9_n136, mult_9_n169);
	or gate_mult_9_n137 (mult_9_n137, mult_9_n135, mult_9_n134);
	xor gate_mult_9_n138 (mult_9_n138, mult_9_n169, mult_9_n136);
	xor gate_mult_9_n131 (mult_9_n131, mult_9_n164, mult_9_n143);
	and gate_mult_9_n130 (mult_9_n130, mult_9_n143, mult_9_n164);
	and gate_mult_9_n129 (mult_9_n129, mult_9_n131, mult_9_n138);
	or gate_mult_9_n132 (mult_9_n132, mult_9_n130, mult_9_n129);
	xor gate_mult_9_n133 (mult_9_n133, mult_9_n138, mult_9_n131);
	xor gate_mult_9_n126 (mult_9_n126, mult_9_n283, mult_9_n276);
	and gate_mult_9_n125 (mult_9_n125, mult_9_n276, mult_9_n283);
	and gate_mult_9_n124 (mult_9_n124, mult_9_n126, mult_9_n269);
	or gate_mult_9_n127 (mult_9_n127, mult_9_n125, mult_9_n124);
	xor gate_mult_9_n128 (mult_9_n128, mult_9_n269, mult_9_n126);
	xor gate_mult_9_n121 (mult_9_n121, mult_9_n262, mult_9_n255);
	and gate_mult_9_n120 (mult_9_n120, mult_9_n255, mult_9_n262);
	and gate_mult_9_n119 (mult_9_n119, mult_9_n121, mult_9_n248);
	or gate_mult_9_n122 (mult_9_n122, mult_9_n120, mult_9_n119);
	xor gate_mult_9_n123 (mult_9_n123, mult_9_n248, mult_9_n121);
	xor gate_mult_9_n116 (mult_9_n116, mult_9_n154, mult_9_n152);
	and gate_mult_9_n115 (mult_9_n115, mult_9_n152, mult_9_n154);
	and gate_mult_9_n114 (mult_9_n114, mult_9_n116, mult_9_n147);
	or gate_mult_9_n117 (mult_9_n117, mult_9_n115, mult_9_n114);
	xor gate_mult_9_n118 (mult_9_n118, mult_9_n147, mult_9_n116);
	xor gate_mult_9_n111 (mult_9_n111, mult_9_n123, mult_9_n128);
	and gate_mult_9_n110 (mult_9_n110, mult_9_n128, mult_9_n123);
	and gate_mult_9_n109 (mult_9_n109, mult_9_n142, mult_9_n111);
	or gate_mult_9_n112 (mult_9_n112, mult_9_n110, mult_9_n109);
	xor gate_mult_9_n113 (mult_9_n113, mult_9_n111, mult_9_n142);
	xor gate_mult_9_n106 (mult_9_n106, mult_9_n118, mult_9_n137);
	and gate_mult_9_n105 (mult_9_n105, mult_9_n137, mult_9_n118);
	and gate_mult_9_n104 (mult_9_n104, mult_9_n106, mult_9_n113);
	or gate_mult_9_n107 (mult_9_n107, mult_9_n105, mult_9_n104);
	xor gate_mult_9_n108 (mult_9_n108, mult_9_n113, mult_9_n106);
	xor gate_mult_9_n101 (mult_9_n101, mult_9_n275, mult_9_n268);
	and gate_mult_9_n100 (mult_9_n100, mult_9_n268, mult_9_n275);
	and gate_mult_9_n99 (mult_9_n99, mult_9_n101, mult_9_n261);
	or gate_mult_9_n102 (mult_9_n102, mult_9_n100, mult_9_n99);
	xor gate_mult_9_n103 (mult_9_n103, mult_9_n261, mult_9_n101);
	xor gate_mult_9_n96 (mult_9_n96, mult_9_n254, mult_9_n247);
	and gate_mult_9_n95 (mult_9_n95, mult_9_n247, mult_9_n254);
	and gate_mult_9_n94 (mult_9_n94, mult_9_n127, mult_9_n96);
	or gate_mult_9_n97 (mult_9_n97, mult_9_n95, mult_9_n94);
	xor gate_mult_9_n98 (mult_9_n98, mult_9_n96, mult_9_n127);
	xor gate_mult_9_n91 (mult_9_n91, mult_9_n122, mult_9_n103);
	and gate_mult_9_n90 (mult_9_n90, mult_9_n103, mult_9_n122);
	and gate_mult_9_n89 (mult_9_n89, mult_9_n91, mult_9_n98);
	or gate_mult_9_n92 (mult_9_n92, mult_9_n90, mult_9_n89);
	xor gate_mult_9_n93 (mult_9_n93, mult_9_n98, mult_9_n91);
	xor gate_mult_9_n86 (mult_9_n86, mult_9_n117, mult_9_n93);
	and gate_mult_9_n85 (mult_9_n85, mult_9_n93, mult_9_n117);
	and gate_mult_9_n84 (mult_9_n84, mult_9_n86, mult_9_n112);
	or gate_mult_9_n87 (mult_9_n87, mult_9_n85, mult_9_n84);
	xor gate_mult_9_n88 (mult_9_n88, mult_9_n112, mult_9_n86);
	xor gate_mult_9_n81 (mult_9_n81, mult_9_n267, mult_9_n260);
	and gate_mult_9_n80 (mult_9_n80, mult_9_n260, mult_9_n267);
	and gate_mult_9_n79 (mult_9_n79, mult_9_n81, mult_9_n253);
	or gate_mult_9_n82 (mult_9_n82, mult_9_n80, mult_9_n79);
	xor gate_mult_9_n83 (mult_9_n83, mult_9_n253, mult_9_n81);
	xor gate_mult_9_n76 (mult_9_n76, mult_9_n246, mult_9_n102);
	and gate_mult_9_n75 (mult_9_n75, mult_9_n102, mult_9_n246);
	and gate_mult_9_n74 (mult_9_n74, mult_9_n76, mult_9_n83);
	or gate_mult_9_n77 (mult_9_n77, mult_9_n75, mult_9_n74);
	xor gate_mult_9_n78 (mult_9_n78, mult_9_n83, mult_9_n76);
	xor gate_mult_9_n71 (mult_9_n71, mult_9_n97, mult_9_n92);
	and gate_mult_9_n70 (mult_9_n70, mult_9_n92, mult_9_n97);
	and gate_mult_9_n69 (mult_9_n69, mult_9_n71, mult_9_n78);
	or gate_mult_9_n72 (mult_9_n72, mult_9_n70, mult_9_n69);
	xor gate_mult_9_n73 (mult_9_n73, mult_9_n78, mult_9_n71);
	xor gate_mult_9_n66 (mult_9_n66, mult_9_n259, mult_9_n252);
	and gate_mult_9_n65 (mult_9_n65, mult_9_n252, mult_9_n259);
	and gate_mult_9_n64 (mult_9_n64, mult_9_n66, mult_9_n245);
	or gate_mult_9_n67 (mult_9_n67, mult_9_n65, mult_9_n64);
	xor gate_mult_9_n68 (mult_9_n68, mult_9_n245, mult_9_n66);
	xor gate_mult_9_n61 (mult_9_n61, mult_9_n82, mult_9_n68);
	and gate_mult_9_n60 (mult_9_n60, mult_9_n68, mult_9_n82);
	and gate_mult_9_n59 (mult_9_n59, mult_9_n77, mult_9_n61);
	or gate_mult_9_n62 (mult_9_n62, mult_9_n60, mult_9_n59);
	xor gate_mult_9_n63 (mult_9_n63, mult_9_n61, mult_9_n77);
	xor gate_mult_9_n56 (mult_9_n56, mult_9_n251, mult_9_n244);
	and gate_mult_9_n55 (mult_9_n55, mult_9_n244, mult_9_n251);
	and gate_mult_9_n54 (mult_9_n54, mult_9_n67, mult_9_n56);
	or gate_mult_9_n57 (mult_9_n57, mult_9_n55, mult_9_n54);
	xor gate_mult_9_n58 (mult_9_n58, mult_9_n56, mult_9_n67);
	and gate_mult_9_n53 (mult_9_n53, mult_9_n305, mult_9_n298);
	xor gate_sum_1 (sum_1, mult_9_n298, mult_9_n305);
	xor gate_mult_9_n39 (mult_9_n39, mult_9_n290, mult_9_n242);
	and gate_mult_9_n38 (mult_9_n38, mult_9_n242, mult_9_n290);
	and gate_mult_9_n37 (mult_9_n37, mult_9_n39, mult_9_n53);
	or gate_mult_9_n52 (mult_9_n52, mult_9_n38, mult_9_n37);
	xor gate_sum_2 (sum_2, mult_9_n53, mult_9_n39);
	xor gate_mult_9_n36 (mult_9_n36, mult_9_n240, mult_9_n238);
	and gate_mult_9_n35 (mult_9_n35, mult_9_n238, mult_9_n240);
	and gate_mult_9_n34 (mult_9_n34, mult_9_n36, mult_9_n52);
	or gate_mult_9_n51 (mult_9_n51, mult_9_n35, mult_9_n34);
	xor gate_sum_3 (sum_3, mult_9_n52, mult_9_n36);
	xor gate_mult_9_n33 (mult_9_n33, mult_9_n231, mult_9_n226);
	and gate_mult_9_n32 (mult_9_n32, mult_9_n226, mult_9_n231);
	and gate_mult_9_n31 (mult_9_n31, mult_9_n33, mult_9_n51);
	or gate_mult_9_n50 (mult_9_n50, mult_9_n32, mult_9_n31);
	xor gate_sum_4 (sum_4, mult_9_n51, mult_9_n33);
	xor gate_mult_9_n30 (mult_9_n30, mult_9_n225, mult_9_n209);
	and gate_mult_9_n29 (mult_9_n29, mult_9_n209, mult_9_n225);
	and gate_mult_9_n28 (mult_9_n28, mult_9_n30, mult_9_n50);
	or gate_mult_9_n49 (mult_9_n49, mult_9_n29, mult_9_n28);
	xor gate_sum_5 (sum_5, mult_9_n50, mult_9_n30);
	xor gate_mult_9_n27 (mult_9_n27, mult_9_n192, mult_9_n187);
	and gate_mult_9_n26 (mult_9_n26, mult_9_n187, mult_9_n192);
	and gate_mult_9_n25 (mult_9_n25, mult_9_n27, mult_9_n49);
	or gate_mult_9_n48 (mult_9_n48, mult_9_n26, mult_9_n25);
	xor gate_sum_6 (sum_6, mult_9_n49, mult_9_n27);
	xor gate_mult_9_n24 (mult_9_n24, mult_9_n186, mult_9_n160);
	and gate_mult_9_n23 (mult_9_n23, mult_9_n160, mult_9_n186);
	and gate_mult_9_n22 (mult_9_n22, mult_9_n48, mult_9_n24);
	or gate_mult_9_n47 (mult_9_n47, mult_9_n23, mult_9_n22);
	xor gate_sum_7 (sum_7, mult_9_n24, mult_9_n48);
	xor gate_mult_9_n21 (mult_9_n21, mult_9_n159, mult_9_n133);
	and gate_mult_9_n20 (mult_9_n20, mult_9_n133, mult_9_n159);
	and gate_mult_9_n19 (mult_9_n19, mult_9_n47, mult_9_n21);
	or gate_mult_9_n46 (mult_9_n46, mult_9_n20, mult_9_n19);
	xor gate_sum_8 (sum_8, mult_9_n21, mult_9_n47);
	xor gate_mult_9_n18 (mult_9_n18, mult_9_n132, mult_9_n108);
	and gate_mult_9_n17 (mult_9_n17, mult_9_n108, mult_9_n132);
	and gate_mult_9_n16 (mult_9_n16, mult_9_n46, mult_9_n18);
	or gate_mult_9_n45 (mult_9_n45, mult_9_n17, mult_9_n16);
	xor gate_sum_9 (sum_9, mult_9_n18, mult_9_n46);
	xor gate_mult_9_n15 (mult_9_n15, mult_9_n107, mult_9_n88);
	and gate_mult_9_n14 (mult_9_n14, mult_9_n88, mult_9_n107);
	and gate_mult_9_n13 (mult_9_n13, mult_9_n45, mult_9_n15);
	or gate_mult_9_n44 (mult_9_n44, mult_9_n14, mult_9_n13);
	xor gate_sum_10 (sum_10, mult_9_n15, mult_9_n45);
	xor gate_mult_9_n12 (mult_9_n12, mult_9_n87, mult_9_n73);
	and gate_mult_9_n11 (mult_9_n11, mult_9_n73, mult_9_n87);
	and gate_mult_9_n10 (mult_9_n10, mult_9_n44, mult_9_n12);
	or gate_mult_9_n43 (mult_9_n43, mult_9_n11, mult_9_n10);
	xor gate_sum_11 (sum_11, mult_9_n12, mult_9_n44);
	xor gate_mult_9_n9 (mult_9_n9, mult_9_n63, mult_9_n72);
	and gate_mult_9_n8 (mult_9_n8, mult_9_n72, mult_9_n63);
	and gate_mult_9_n7 (mult_9_n7, mult_9_n43, mult_9_n9);
	or gate_mult_9_n42 (mult_9_n42, mult_9_n8, mult_9_n7);
	xor gate_sum_12 (sum_12, mult_9_n9, mult_9_n43);
	xor gate_mult_9_n6 (mult_9_n6, mult_9_n58, mult_9_n62);
	and gate_mult_9_n5 (mult_9_n5, mult_9_n62, mult_9_n58);
	and gate_mult_9_n4 (mult_9_n4, mult_9_n42, mult_9_n6);
	or gate_mult_9_n41 (mult_9_n41, mult_9_n5, mult_9_n4);
	xor gate_sum_13 (sum_13, mult_9_n6, mult_9_n42);
	xor gate_mult_9_n3 (mult_9_n3, mult_9_n243, mult_9_n57);
	and gate_mult_9_n2 (mult_9_n2, mult_9_n57, mult_9_n243);
	and gate_mult_9_n1 (mult_9_n1, mult_9_n41, mult_9_n3);
	or gate_mult_9_n40 (mult_9_n40, mult_9_n2, mult_9_n1);
	xor gate_sum_14 (sum_14, mult_9_n3, mult_9_n41);
	buf gate_sum_15 (sum_15, mult_9_n40);
endmodule

