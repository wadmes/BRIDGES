
module test (a_0, a_1, a_2, a_3, a_4, a_5, a_6, a_7, a_8, a_9, a_10, a_11, a_12, a_13, a_14, a_15, 
   b_0, b_1, b_2, b_3, b_4, b_5, b_6, b_7, b_8, b_9, b_10, b_11, b_12, b_13, b_14, b_15,
   sum_0, sum_1, sum_2, sum_3, sum_4, sum_5, sum_6, sum_7, sum_8, sum_9, sum_10, sum_11, 
   sum_12, sum_13, sum_14, sum_15, sum_16, sum_17, sum_18, sum_19, sum_20, sum_21, sum_22, 
   sum_23, sum_24, sum_25, sum_26, sum_27, sum_28, sum_29, sum_30, sum_31);

  input a_0;
  input a_1;
  input a_2;
  input a_3;
  input a_4;
  input a_5;
  input a_6;
  input a_7;
  input a_8;
  input a_9;
  input a_10;
  input a_11;
  input a_12;
  input a_13;
  input a_14;
  input a_15;

  input b_0;
  input b_1;
  input b_2;
  input b_3;
  input b_4;
  input b_5;
  input b_6;
  input b_7;
  input b_8;
  input b_9;
  input b_10;
  input b_11;
  input b_12;
  input b_13;
  input b_14;
  input b_15;


  output sum_0;
  output sum_1;
  output sum_2;
  output sum_3;
  output sum_4;
  output sum_5;
  output sum_6;
  output sum_7;
  output sum_8;
  output sum_9;
  output sum_10;
  output sum_11;
  output sum_12;
  output sum_13;
  output sum_14;
  output sum_15;
  output sum_16;
output sum_17;
output sum_18;
output sum_19;
output sum_20;
output sum_21;
output sum_22;
output sum_23;
output sum_24;
output sum_25;
output sum_26;
output sum_27;
output sum_28;
output sum_29;
output sum_30;
output sum_31;
  

	not gate_anoymous_9_n1403 (anoymous_9_n1403, a_0);
	xor gate_anoymous_9_n1386 (anoymous_9_n1386, a_1, a_0);
	nand gate_anoymous_9_n1394 (anoymous_9_n1394, anoymous_9_n1403, anoymous_9_n1386);
	xnor gate_anoymous_9_n1402 (anoymous_9_n1402, a_1, a_2);
	xor gate_anoymous_9_n1385 (anoymous_9_n1385, a_3, a_2);
	nand gate_anoymous_9_n1393 (anoymous_9_n1393, anoymous_9_n1385, anoymous_9_n1402);
	xnor gate_anoymous_9_n1401 (anoymous_9_n1401, a_3, a_4);
	xor gate_anoymous_9_n1384 (anoymous_9_n1384, a_5, a_4);
	nand gate_anoymous_9_n1392 (anoymous_9_n1392, anoymous_9_n1384, anoymous_9_n1401);
	xnor gate_anoymous_9_n1400 (anoymous_9_n1400, a_5, a_6);
	xor gate_anoymous_9_n1383 (anoymous_9_n1383, a_7, a_6);
	nand gate_anoymous_9_n1391 (anoymous_9_n1391, anoymous_9_n1383, anoymous_9_n1400);
	xnor gate_anoymous_9_n1399 (anoymous_9_n1399, a_7, a_8);
	xor gate_anoymous_9_n1382 (anoymous_9_n1382, a_9, a_8);
	nand gate_anoymous_9_n1390 (anoymous_9_n1390, anoymous_9_n1382, anoymous_9_n1399);
	xnor gate_anoymous_9_n1398 (anoymous_9_n1398, a_9, a_10);
	xor gate_anoymous_9_n1381 (anoymous_9_n1381, a_11, a_10);
	nand gate_anoymous_9_n1389 (anoymous_9_n1389, anoymous_9_n1381, anoymous_9_n1398);
	xnor gate_anoymous_9_n1397 (anoymous_9_n1397, a_11, a_12);
	xor gate_anoymous_9_n1380 (anoymous_9_n1380, a_13, a_12);
	nand gate_anoymous_9_n1388 (anoymous_9_n1388, anoymous_9_n1380, anoymous_9_n1397);
	xnor gate_anoymous_9_n1396 (anoymous_9_n1396, a_13, a_14);
	xor gate_anoymous_9_n1379 (anoymous_9_n1379, a_15, a_14);
	nand gate_anoymous_9_n1387 (anoymous_9_n1387, anoymous_9_n1379, anoymous_9_n1396);
	not gate_anoymous_9_n1420 (anoymous_9_n1420, a_15);
	not gate_anoymous_9_n1411 (anoymous_9_n1411, anoymous_9_n1);
	not gate_anoymous_9_n1410 (anoymous_9_n1410, anoymous_9_n7);
	not gate_anoymous_9_n1409 (anoymous_9_n1409, anoymous_9_n13);
	not gate_anoymous_9_n1408 (anoymous_9_n1408, anoymous_9_n19);
	not gate_anoymous_9_n1407 (anoymous_9_n1407, anoymous_9_n25);
	not gate_anoymous_9_n1406 (anoymous_9_n1406, anoymous_9_n31);
	not gate_anoymous_9_n1405 (anoymous_9_n1405, anoymous_9_n37);
	not gate_anoymous_9_n1404 (anoymous_9_n1404, anoymous_9_n43);
	buf gate_anoymous_9_n1395 (anoymous_9_n1395, anoymous_9_n1420);
	buf gate_anoymous_9_n1377 (anoymous_9_n1377, b_1);
	buf gate_anoymous_9_n1376 (anoymous_9_n1376, b_2);
	buf gate_anoymous_9_n1375 (anoymous_9_n1375, b_3);
	buf gate_anoymous_9_n1374 (anoymous_9_n1374, b_4);
	buf gate_anoymous_9_n1373 (anoymous_9_n1373, b_5);
	buf gate_anoymous_9_n1372 (anoymous_9_n1372, b_6);
	buf gate_anoymous_9_n1371 (anoymous_9_n1371, b_7);
	buf gate_anoymous_9_n1370 (anoymous_9_n1370, b_8);
	buf gate_anoymous_9_n1369 (anoymous_9_n1369, b_9);
	buf gate_anoymous_9_n1368 (anoymous_9_n1368, b_10);
	buf gate_anoymous_9_n1367 (anoymous_9_n1367, b_11);
	buf gate_anoymous_9_n1366 (anoymous_9_n1366, b_12);
	buf gate_anoymous_9_n1365 (anoymous_9_n1365, b_13);
	buf gate_anoymous_9_n1364 (anoymous_9_n1364, b_14);
	buf gate_anoymous_9_n1363 (anoymous_9_n1363, b_15);
	or gate_anoymous_9_n1362 (anoymous_9_n1362, anoymous_9_n49, anoymous_9_n1411);
	xnor gate_anoymous_9_n1361 (anoymous_9_n1361, anoymous_9_n49, anoymous_9_n1);
	xnor gate_anoymous_9_n1360 (anoymous_9_n1360, anoymous_9_n1377, anoymous_9_n1);
	xnor gate_anoymous_9_n1359 (anoymous_9_n1359, anoymous_9_n1376, anoymous_9_n1);
	xnor gate_anoymous_9_n1358 (anoymous_9_n1358, anoymous_9_n1375, anoymous_9_n1);
	xnor gate_anoymous_9_n1357 (anoymous_9_n1357, anoymous_9_n1374, anoymous_9_n1);
	xnor gate_anoymous_9_n1356 (anoymous_9_n1356, anoymous_9_n1373, anoymous_9_n1);
	xnor gate_anoymous_9_n1355 (anoymous_9_n1355, anoymous_9_n1372, anoymous_9_n1);
	xnor gate_anoymous_9_n1354 (anoymous_9_n1354, anoymous_9_n1371, anoymous_9_n1);
	xnor gate_anoymous_9_n1353 (anoymous_9_n1353, anoymous_9_n1370, anoymous_9_n1);
	xnor gate_anoymous_9_n1352 (anoymous_9_n1352, anoymous_9_n1369, anoymous_9_n1);
	xnor gate_anoymous_9_n1351 (anoymous_9_n1351, anoymous_9_n1368, anoymous_9_n1);
	xnor gate_anoymous_9_n1350 (anoymous_9_n1350, anoymous_9_n1367, anoymous_9_n1);
	xnor gate_anoymous_9_n1349 (anoymous_9_n1349, anoymous_9_n1366, anoymous_9_n1);
	xnor gate_anoymous_9_n1348 (anoymous_9_n1348, anoymous_9_n1365, anoymous_9_n1);
	xnor gate_anoymous_9_n1347 (anoymous_9_n1347, anoymous_9_n1364, anoymous_9_n1);
	xnor gate_anoymous_9_n1346 (anoymous_9_n1346, anoymous_9_n1363, anoymous_9_n1);
	not gate_anoymous_9_n1050 (anoymous_9_n1050, anoymous_9_n3);
	and gate_sum_0 (sum_0, anoymous_9_n49, anoymous_9_n1050);
	or gate_anoymous_9_n1049 (anoymous_9_n1049, anoymous_9_n5, anoymous_9_n1361);
	or gate_anoymous_9_n1048 (anoymous_9_n1048, anoymous_9_n1360, anoymous_9_n3);
	nand gate_anoymous_9_n1211 (anoymous_9_n1211, anoymous_9_n1049, anoymous_9_n1048);
	or gate_anoymous_9_n1047 (anoymous_9_n1047, anoymous_9_n5, anoymous_9_n1360);
	or gate_anoymous_9_n1046 (anoymous_9_n1046, anoymous_9_n1359, anoymous_9_n3);
	nand gate_anoymous_9_n1210 (anoymous_9_n1210, anoymous_9_n1047, anoymous_9_n1046);
	or gate_anoymous_9_n1045 (anoymous_9_n1045, anoymous_9_n5, anoymous_9_n1359);
	or gate_anoymous_9_n1044 (anoymous_9_n1044, anoymous_9_n1358, anoymous_9_n3);
	nand gate_anoymous_9_n1209 (anoymous_9_n1209, anoymous_9_n1045, anoymous_9_n1044);
	or gate_anoymous_9_n1043 (anoymous_9_n1043, anoymous_9_n5, anoymous_9_n1358);
	or gate_anoymous_9_n1042 (anoymous_9_n1042, anoymous_9_n1357, anoymous_9_n3);
	nand gate_anoymous_9_n1208 (anoymous_9_n1208, anoymous_9_n1043, anoymous_9_n1042);
	or gate_anoymous_9_n1041 (anoymous_9_n1041, anoymous_9_n5, anoymous_9_n1357);
	or gate_anoymous_9_n1040 (anoymous_9_n1040, anoymous_9_n1356, anoymous_9_n3);
	nand gate_anoymous_9_n1207 (anoymous_9_n1207, anoymous_9_n1041, anoymous_9_n1040);
	or gate_anoymous_9_n1039 (anoymous_9_n1039, anoymous_9_n5, anoymous_9_n1356);
	or gate_anoymous_9_n1038 (anoymous_9_n1038, anoymous_9_n1355, anoymous_9_n3);
	nand gate_anoymous_9_n1206 (anoymous_9_n1206, anoymous_9_n1039, anoymous_9_n1038);
	or gate_anoymous_9_n1037 (anoymous_9_n1037, anoymous_9_n5, anoymous_9_n1355);
	or gate_anoymous_9_n1036 (anoymous_9_n1036, anoymous_9_n1354, anoymous_9_n3);
	nand gate_anoymous_9_n1205 (anoymous_9_n1205, anoymous_9_n1037, anoymous_9_n1036);
	or gate_anoymous_9_n1035 (anoymous_9_n1035, anoymous_9_n5, anoymous_9_n1354);
	or gate_anoymous_9_n1034 (anoymous_9_n1034, anoymous_9_n1353, anoymous_9_n3);
	nand gate_anoymous_9_n1204 (anoymous_9_n1204, anoymous_9_n1035, anoymous_9_n1034);
	or gate_anoymous_9_n1033 (anoymous_9_n1033, anoymous_9_n5, anoymous_9_n1353);
	or gate_anoymous_9_n1032 (anoymous_9_n1032, anoymous_9_n1352, anoymous_9_n4);
	nand gate_anoymous_9_n1203 (anoymous_9_n1203, anoymous_9_n1033, anoymous_9_n1032);
	or gate_anoymous_9_n1031 (anoymous_9_n1031, anoymous_9_n6, anoymous_9_n1352);
	or gate_anoymous_9_n1030 (anoymous_9_n1030, anoymous_9_n1351, anoymous_9_n4);
	nand gate_anoymous_9_n1202 (anoymous_9_n1202, anoymous_9_n1031, anoymous_9_n1030);
	or gate_anoymous_9_n1029 (anoymous_9_n1029, anoymous_9_n6, anoymous_9_n1351);
	or gate_anoymous_9_n1028 (anoymous_9_n1028, anoymous_9_n1350, anoymous_9_n4);
	nand gate_anoymous_9_n1201 (anoymous_9_n1201, anoymous_9_n1029, anoymous_9_n1028);
	or gate_anoymous_9_n1027 (anoymous_9_n1027, anoymous_9_n6, anoymous_9_n1350);
	or gate_anoymous_9_n1026 (anoymous_9_n1026, anoymous_9_n1349, anoymous_9_n4);
	nand gate_anoymous_9_n1200 (anoymous_9_n1200, anoymous_9_n1027, anoymous_9_n1026);
	or gate_anoymous_9_n1025 (anoymous_9_n1025, anoymous_9_n6, anoymous_9_n1349);
	or gate_anoymous_9_n1024 (anoymous_9_n1024, anoymous_9_n1348, anoymous_9_n4);
	nand gate_anoymous_9_n1199 (anoymous_9_n1199, anoymous_9_n1025, anoymous_9_n1024);
	or gate_anoymous_9_n1023 (anoymous_9_n1023, anoymous_9_n6, anoymous_9_n1348);
	or gate_anoymous_9_n1022 (anoymous_9_n1022, anoymous_9_n1347, anoymous_9_n4);
	nand gate_anoymous_9_n1198 (anoymous_9_n1198, anoymous_9_n1023, anoymous_9_n1022);
	or gate_anoymous_9_n1021 (anoymous_9_n1021, anoymous_9_n6, anoymous_9_n1347);
	or gate_anoymous_9_n1020 (anoymous_9_n1020, anoymous_9_n1346, anoymous_9_n4);
	nand gate_anoymous_9_n1197 (anoymous_9_n1197, anoymous_9_n1021, anoymous_9_n1020);
	or gate_anoymous_9_n1019 (anoymous_9_n1019, anoymous_9_n6, anoymous_9_n1346);
	or gate_anoymous_9_n1018 (anoymous_9_n1018, anoymous_9_n1411, anoymous_9_n4);
	nand gate_anoymous_9_n1196 (anoymous_9_n1196, anoymous_9_n1019, anoymous_9_n1018);
	and gate_anoymous_9_n1017 (anoymous_9_n1017, anoymous_9_n6, anoymous_9_n4);
	or gate_anoymous_9_n1195 (anoymous_9_n1195, anoymous_9_n1411, anoymous_9_n1017);
	or gate_anoymous_9_n1016 (anoymous_9_n1016, anoymous_9_n1362, anoymous_9_n4);
	or gate_anoymous_9_n1015 (anoymous_9_n1015, anoymous_9_n6, anoymous_9_n1411);
	nand gate_anoymous_9_n1059 (anoymous_9_n1059, anoymous_9_n1016, anoymous_9_n1015);
	or gate_anoymous_9_n1345 (anoymous_9_n1345, anoymous_9_n49, anoymous_9_n1410);
	xnor gate_anoymous_9_n1344 (anoymous_9_n1344, anoymous_9_n49, anoymous_9_n7);
	xnor gate_anoymous_9_n1343 (anoymous_9_n1343, anoymous_9_n1377, anoymous_9_n7);
	xnor gate_anoymous_9_n1342 (anoymous_9_n1342, anoymous_9_n1376, anoymous_9_n7);
	xnor gate_anoymous_9_n1341 (anoymous_9_n1341, anoymous_9_n1375, anoymous_9_n7);
	xnor gate_anoymous_9_n1340 (anoymous_9_n1340, anoymous_9_n1374, anoymous_9_n7);
	xnor gate_anoymous_9_n1339 (anoymous_9_n1339, anoymous_9_n1373, anoymous_9_n7);
	xnor gate_anoymous_9_n1338 (anoymous_9_n1338, anoymous_9_n1372, anoymous_9_n7);
	xnor gate_anoymous_9_n1337 (anoymous_9_n1337, anoymous_9_n1371, anoymous_9_n7);
	xnor gate_anoymous_9_n1336 (anoymous_9_n1336, anoymous_9_n1370, anoymous_9_n7);
	xnor gate_anoymous_9_n1335 (anoymous_9_n1335, anoymous_9_n1369, anoymous_9_n7);
	xnor gate_anoymous_9_n1334 (anoymous_9_n1334, anoymous_9_n1368, anoymous_9_n7);
	xnor gate_anoymous_9_n1333 (anoymous_9_n1333, anoymous_9_n1367, anoymous_9_n7);
	xnor gate_anoymous_9_n1332 (anoymous_9_n1332, anoymous_9_n1366, anoymous_9_n7);
	xnor gate_anoymous_9_n1331 (anoymous_9_n1331, anoymous_9_n1365, anoymous_9_n7);
	xnor gate_anoymous_9_n1330 (anoymous_9_n1330, anoymous_9_n1364, anoymous_9_n7);
	xnor gate_anoymous_9_n1329 (anoymous_9_n1329, anoymous_9_n1363, anoymous_9_n7);
	not gate_anoymous_9_n1013 (anoymous_9_n1013, anoymous_9_n9);
	and gate_anoymous_9_n1194 (anoymous_9_n1194, anoymous_9_n49, anoymous_9_n1013);
	or gate_anoymous_9_n1012 (anoymous_9_n1012, anoymous_9_n11, anoymous_9_n1344);
	or gate_anoymous_9_n1011 (anoymous_9_n1011, anoymous_9_n9, anoymous_9_n1343);
	nand gate_anoymous_9_n1193 (anoymous_9_n1193, anoymous_9_n1012, anoymous_9_n1011);
	or gate_anoymous_9_n1010 (anoymous_9_n1010, anoymous_9_n11, anoymous_9_n1343);
	or gate_anoymous_9_n1009 (anoymous_9_n1009, anoymous_9_n9, anoymous_9_n1342);
	nand gate_anoymous_9_n1192 (anoymous_9_n1192, anoymous_9_n1010, anoymous_9_n1009);
	or gate_anoymous_9_n1008 (anoymous_9_n1008, anoymous_9_n11, anoymous_9_n1342);
	or gate_anoymous_9_n1007 (anoymous_9_n1007, anoymous_9_n9, anoymous_9_n1341);
	nand gate_anoymous_9_n1191 (anoymous_9_n1191, anoymous_9_n1008, anoymous_9_n1007);
	or gate_anoymous_9_n1006 (anoymous_9_n1006, anoymous_9_n11, anoymous_9_n1341);
	or gate_anoymous_9_n1005 (anoymous_9_n1005, anoymous_9_n9, anoymous_9_n1340);
	nand gate_anoymous_9_n1190 (anoymous_9_n1190, anoymous_9_n1006, anoymous_9_n1005);
	or gate_anoymous_9_n1004 (anoymous_9_n1004, anoymous_9_n11, anoymous_9_n1340);
	or gate_anoymous_9_n1003 (anoymous_9_n1003, anoymous_9_n9, anoymous_9_n1339);
	nand gate_anoymous_9_n1189 (anoymous_9_n1189, anoymous_9_n1004, anoymous_9_n1003);
	or gate_anoymous_9_n1002 (anoymous_9_n1002, anoymous_9_n11, anoymous_9_n1339);
	or gate_anoymous_9_n1001 (anoymous_9_n1001, anoymous_9_n9, anoymous_9_n1338);
	nand gate_anoymous_9_n1188 (anoymous_9_n1188, anoymous_9_n1002, anoymous_9_n1001);
	or gate_anoymous_9_n1000 (anoymous_9_n1000, anoymous_9_n11, anoymous_9_n1338);
	or gate_anoymous_9_n999 (anoymous_9_n999, anoymous_9_n9, anoymous_9_n1337);
	nand gate_anoymous_9_n1187 (anoymous_9_n1187, anoymous_9_n1000, anoymous_9_n999);
	or gate_anoymous_9_n998 (anoymous_9_n998, anoymous_9_n11, anoymous_9_n1337);
	or gate_anoymous_9_n997 (anoymous_9_n997, anoymous_9_n9, anoymous_9_n1336);
	nand gate_anoymous_9_n1186 (anoymous_9_n1186, anoymous_9_n998, anoymous_9_n997);
	or gate_anoymous_9_n996 (anoymous_9_n996, anoymous_9_n11, anoymous_9_n1336);
	or gate_anoymous_9_n995 (anoymous_9_n995, anoymous_9_n10, anoymous_9_n1335);
	nand gate_anoymous_9_n1185 (anoymous_9_n1185, anoymous_9_n996, anoymous_9_n995);
	or gate_anoymous_9_n994 (anoymous_9_n994, anoymous_9_n12, anoymous_9_n1335);
	or gate_anoymous_9_n993 (anoymous_9_n993, anoymous_9_n10, anoymous_9_n1334);
	nand gate_anoymous_9_n1184 (anoymous_9_n1184, anoymous_9_n994, anoymous_9_n993);
	or gate_anoymous_9_n992 (anoymous_9_n992, anoymous_9_n12, anoymous_9_n1334);
	or gate_anoymous_9_n991 (anoymous_9_n991, anoymous_9_n10, anoymous_9_n1333);
	nand gate_anoymous_9_n1183 (anoymous_9_n1183, anoymous_9_n992, anoymous_9_n991);
	or gate_anoymous_9_n990 (anoymous_9_n990, anoymous_9_n12, anoymous_9_n1333);
	or gate_anoymous_9_n989 (anoymous_9_n989, anoymous_9_n10, anoymous_9_n1332);
	nand gate_anoymous_9_n1182 (anoymous_9_n1182, anoymous_9_n990, anoymous_9_n989);
	or gate_anoymous_9_n988 (anoymous_9_n988, anoymous_9_n12, anoymous_9_n1332);
	or gate_anoymous_9_n987 (anoymous_9_n987, anoymous_9_n10, anoymous_9_n1331);
	nand gate_anoymous_9_n1181 (anoymous_9_n1181, anoymous_9_n988, anoymous_9_n987);
	or gate_anoymous_9_n986 (anoymous_9_n986, anoymous_9_n12, anoymous_9_n1331);
	or gate_anoymous_9_n985 (anoymous_9_n985, anoymous_9_n10, anoymous_9_n1330);
	nand gate_anoymous_9_n1180 (anoymous_9_n1180, anoymous_9_n986, anoymous_9_n985);
	or gate_anoymous_9_n984 (anoymous_9_n984, anoymous_9_n12, anoymous_9_n1330);
	or gate_anoymous_9_n983 (anoymous_9_n983, anoymous_9_n10, anoymous_9_n1329);
	nand gate_anoymous_9_n1179 (anoymous_9_n1179, anoymous_9_n984, anoymous_9_n983);
	or gate_anoymous_9_n982 (anoymous_9_n982, anoymous_9_n12, anoymous_9_n1329);
	or gate_anoymous_9_n981 (anoymous_9_n981, anoymous_9_n10, anoymous_9_n1410);
	nand gate_anoymous_9_n1178 (anoymous_9_n1178, anoymous_9_n982, anoymous_9_n981);
	and gate_anoymous_9_n980 (anoymous_9_n980, anoymous_9_n12, anoymous_9_n10);
	or gate_anoymous_9_n1177 (anoymous_9_n1177, anoymous_9_n1410, anoymous_9_n980);
	or gate_anoymous_9_n979 (anoymous_9_n979, anoymous_9_n10, anoymous_9_n1345);
	or gate_anoymous_9_n978 (anoymous_9_n978, anoymous_9_n12, anoymous_9_n1410);
	nand gate_anoymous_9_n1058 (anoymous_9_n1058, anoymous_9_n979, anoymous_9_n978);
	or gate_anoymous_9_n1328 (anoymous_9_n1328, anoymous_9_n49, anoymous_9_n1409);
	xnor gate_anoymous_9_n1327 (anoymous_9_n1327, anoymous_9_n49, anoymous_9_n13);
	xnor gate_anoymous_9_n1326 (anoymous_9_n1326, anoymous_9_n1377, anoymous_9_n13);
	xnor gate_anoymous_9_n1325 (anoymous_9_n1325, anoymous_9_n1376, anoymous_9_n13);
	xnor gate_anoymous_9_n1324 (anoymous_9_n1324, anoymous_9_n1375, anoymous_9_n13);
	xnor gate_anoymous_9_n1323 (anoymous_9_n1323, anoymous_9_n1374, anoymous_9_n13);
	xnor gate_anoymous_9_n1322 (anoymous_9_n1322, anoymous_9_n1373, anoymous_9_n13);
	xnor gate_anoymous_9_n1321 (anoymous_9_n1321, anoymous_9_n1372, anoymous_9_n13);
	xnor gate_anoymous_9_n1320 (anoymous_9_n1320, anoymous_9_n1371, anoymous_9_n13);
	xnor gate_anoymous_9_n1319 (anoymous_9_n1319, anoymous_9_n1370, anoymous_9_n13);
	xnor gate_anoymous_9_n1318 (anoymous_9_n1318, anoymous_9_n1369, anoymous_9_n13);
	xnor gate_anoymous_9_n1317 (anoymous_9_n1317, anoymous_9_n1368, anoymous_9_n13);
	xnor gate_anoymous_9_n1316 (anoymous_9_n1316, anoymous_9_n1367, anoymous_9_n13);
	xnor gate_anoymous_9_n1315 (anoymous_9_n1315, anoymous_9_n1366, anoymous_9_n13);
	xnor gate_anoymous_9_n1314 (anoymous_9_n1314, anoymous_9_n1365, anoymous_9_n13);
	xnor gate_anoymous_9_n1313 (anoymous_9_n1313, anoymous_9_n1364, anoymous_9_n13);
	xnor gate_anoymous_9_n1312 (anoymous_9_n1312, anoymous_9_n1363, anoymous_9_n13);
	not gate_anoymous_9_n976 (anoymous_9_n976, anoymous_9_n15);
	and gate_anoymous_9_n1176 (anoymous_9_n1176, anoymous_9_n49, anoymous_9_n976);
	or gate_anoymous_9_n975 (anoymous_9_n975, anoymous_9_n17, anoymous_9_n1327);
	or gate_anoymous_9_n974 (anoymous_9_n974, anoymous_9_n15, anoymous_9_n1326);
	nand gate_anoymous_9_n1175 (anoymous_9_n1175, anoymous_9_n975, anoymous_9_n974);
	or gate_anoymous_9_n973 (anoymous_9_n973, anoymous_9_n17, anoymous_9_n1326);
	or gate_anoymous_9_n972 (anoymous_9_n972, anoymous_9_n15, anoymous_9_n1325);
	nand gate_anoymous_9_n1174 (anoymous_9_n1174, anoymous_9_n973, anoymous_9_n972);
	or gate_anoymous_9_n971 (anoymous_9_n971, anoymous_9_n17, anoymous_9_n1325);
	or gate_anoymous_9_n970 (anoymous_9_n970, anoymous_9_n15, anoymous_9_n1324);
	nand gate_anoymous_9_n1173 (anoymous_9_n1173, anoymous_9_n971, anoymous_9_n970);
	or gate_anoymous_9_n969 (anoymous_9_n969, anoymous_9_n17, anoymous_9_n1324);
	or gate_anoymous_9_n968 (anoymous_9_n968, anoymous_9_n15, anoymous_9_n1323);
	nand gate_anoymous_9_n1172 (anoymous_9_n1172, anoymous_9_n969, anoymous_9_n968);
	or gate_anoymous_9_n967 (anoymous_9_n967, anoymous_9_n17, anoymous_9_n1323);
	or gate_anoymous_9_n966 (anoymous_9_n966, anoymous_9_n15, anoymous_9_n1322);
	nand gate_anoymous_9_n1171 (anoymous_9_n1171, anoymous_9_n967, anoymous_9_n966);
	or gate_anoymous_9_n965 (anoymous_9_n965, anoymous_9_n17, anoymous_9_n1322);
	or gate_anoymous_9_n964 (anoymous_9_n964, anoymous_9_n15, anoymous_9_n1321);
	nand gate_anoymous_9_n1170 (anoymous_9_n1170, anoymous_9_n965, anoymous_9_n964);
	or gate_anoymous_9_n963 (anoymous_9_n963, anoymous_9_n17, anoymous_9_n1321);
	or gate_anoymous_9_n962 (anoymous_9_n962, anoymous_9_n15, anoymous_9_n1320);
	nand gate_anoymous_9_n1169 (anoymous_9_n1169, anoymous_9_n963, anoymous_9_n962);
	or gate_anoymous_9_n961 (anoymous_9_n961, anoymous_9_n17, anoymous_9_n1320);
	or gate_anoymous_9_n960 (anoymous_9_n960, anoymous_9_n15, anoymous_9_n1319);
	nand gate_anoymous_9_n1168 (anoymous_9_n1168, anoymous_9_n961, anoymous_9_n960);
	or gate_anoymous_9_n959 (anoymous_9_n959, anoymous_9_n17, anoymous_9_n1319);
	or gate_anoymous_9_n958 (anoymous_9_n958, anoymous_9_n16, anoymous_9_n1318);
	nand gate_anoymous_9_n1167 (anoymous_9_n1167, anoymous_9_n959, anoymous_9_n958);
	or gate_anoymous_9_n957 (anoymous_9_n957, anoymous_9_n18, anoymous_9_n1318);
	or gate_anoymous_9_n956 (anoymous_9_n956, anoymous_9_n16, anoymous_9_n1317);
	nand gate_anoymous_9_n1166 (anoymous_9_n1166, anoymous_9_n957, anoymous_9_n956);
	or gate_anoymous_9_n955 (anoymous_9_n955, anoymous_9_n18, anoymous_9_n1317);
	or gate_anoymous_9_n954 (anoymous_9_n954, anoymous_9_n16, anoymous_9_n1316);
	nand gate_anoymous_9_n1165 (anoymous_9_n1165, anoymous_9_n955, anoymous_9_n954);
	or gate_anoymous_9_n953 (anoymous_9_n953, anoymous_9_n18, anoymous_9_n1316);
	or gate_anoymous_9_n952 (anoymous_9_n952, anoymous_9_n16, anoymous_9_n1315);
	nand gate_anoymous_9_n1164 (anoymous_9_n1164, anoymous_9_n953, anoymous_9_n952);
	or gate_anoymous_9_n951 (anoymous_9_n951, anoymous_9_n18, anoymous_9_n1315);
	or gate_anoymous_9_n950 (anoymous_9_n950, anoymous_9_n16, anoymous_9_n1314);
	nand gate_anoymous_9_n1163 (anoymous_9_n1163, anoymous_9_n951, anoymous_9_n950);
	or gate_anoymous_9_n949 (anoymous_9_n949, anoymous_9_n18, anoymous_9_n1314);
	or gate_anoymous_9_n948 (anoymous_9_n948, anoymous_9_n16, anoymous_9_n1313);
	nand gate_anoymous_9_n1162 (anoymous_9_n1162, anoymous_9_n949, anoymous_9_n948);
	or gate_anoymous_9_n947 (anoymous_9_n947, anoymous_9_n18, anoymous_9_n1313);
	or gate_anoymous_9_n946 (anoymous_9_n946, anoymous_9_n16, anoymous_9_n1312);
	nand gate_anoymous_9_n1161 (anoymous_9_n1161, anoymous_9_n947, anoymous_9_n946);
	or gate_anoymous_9_n945 (anoymous_9_n945, anoymous_9_n18, anoymous_9_n1312);
	or gate_anoymous_9_n944 (anoymous_9_n944, anoymous_9_n16, anoymous_9_n1409);
	nand gate_anoymous_9_n1160 (anoymous_9_n1160, anoymous_9_n945, anoymous_9_n944);
	and gate_anoymous_9_n943 (anoymous_9_n943, anoymous_9_n18, anoymous_9_n16);
	or gate_anoymous_9_n1159 (anoymous_9_n1159, anoymous_9_n1409, anoymous_9_n943);
	or gate_anoymous_9_n942 (anoymous_9_n942, anoymous_9_n16, anoymous_9_n1328);
	or gate_anoymous_9_n941 (anoymous_9_n941, anoymous_9_n18, anoymous_9_n1409);
	nand gate_anoymous_9_n1057 (anoymous_9_n1057, anoymous_9_n942, anoymous_9_n941);
	or gate_anoymous_9_n1311 (anoymous_9_n1311, anoymous_9_n49, anoymous_9_n1408);
	xnor gate_anoymous_9_n1310 (anoymous_9_n1310, anoymous_9_n49, anoymous_9_n19);
	xnor gate_anoymous_9_n1309 (anoymous_9_n1309, anoymous_9_n1377, anoymous_9_n19);
	xnor gate_anoymous_9_n1308 (anoymous_9_n1308, anoymous_9_n1376, anoymous_9_n19);
	xnor gate_anoymous_9_n1307 (anoymous_9_n1307, anoymous_9_n1375, anoymous_9_n19);
	xnor gate_anoymous_9_n1306 (anoymous_9_n1306, anoymous_9_n1374, anoymous_9_n19);
	xnor gate_anoymous_9_n1305 (anoymous_9_n1305, anoymous_9_n1373, anoymous_9_n19);
	xnor gate_anoymous_9_n1304 (anoymous_9_n1304, anoymous_9_n1372, anoymous_9_n19);
	xnor gate_anoymous_9_n1303 (anoymous_9_n1303, anoymous_9_n1371, anoymous_9_n19);
	xnor gate_anoymous_9_n1302 (anoymous_9_n1302, anoymous_9_n1370, anoymous_9_n19);
	xnor gate_anoymous_9_n1301 (anoymous_9_n1301, anoymous_9_n1369, anoymous_9_n19);
	xnor gate_anoymous_9_n1300 (anoymous_9_n1300, anoymous_9_n1368, anoymous_9_n19);
	xnor gate_anoymous_9_n1299 (anoymous_9_n1299, anoymous_9_n1367, anoymous_9_n19);
	xnor gate_anoymous_9_n1298 (anoymous_9_n1298, anoymous_9_n1366, anoymous_9_n19);
	xnor gate_anoymous_9_n1297 (anoymous_9_n1297, anoymous_9_n1365, anoymous_9_n19);
	xnor gate_anoymous_9_n1296 (anoymous_9_n1296, anoymous_9_n1364, anoymous_9_n19);
	xnor gate_anoymous_9_n1295 (anoymous_9_n1295, anoymous_9_n1363, anoymous_9_n19);
	not gate_anoymous_9_n939 (anoymous_9_n939, anoymous_9_n21);
	and gate_anoymous_9_n1158 (anoymous_9_n1158, anoymous_9_n49, anoymous_9_n939);
	or gate_anoymous_9_n938 (anoymous_9_n938, anoymous_9_n23, anoymous_9_n1310);
	or gate_anoymous_9_n937 (anoymous_9_n937, anoymous_9_n21, anoymous_9_n1309);
	nand gate_anoymous_9_n1157 (anoymous_9_n1157, anoymous_9_n938, anoymous_9_n937);
	or gate_anoymous_9_n936 (anoymous_9_n936, anoymous_9_n23, anoymous_9_n1309);
	or gate_anoymous_9_n935 (anoymous_9_n935, anoymous_9_n21, anoymous_9_n1308);
	nand gate_anoymous_9_n1156 (anoymous_9_n1156, anoymous_9_n936, anoymous_9_n935);
	or gate_anoymous_9_n934 (anoymous_9_n934, anoymous_9_n23, anoymous_9_n1308);
	or gate_anoymous_9_n933 (anoymous_9_n933, anoymous_9_n21, anoymous_9_n1307);
	nand gate_anoymous_9_n1155 (anoymous_9_n1155, anoymous_9_n934, anoymous_9_n933);
	or gate_anoymous_9_n932 (anoymous_9_n932, anoymous_9_n23, anoymous_9_n1307);
	or gate_anoymous_9_n931 (anoymous_9_n931, anoymous_9_n21, anoymous_9_n1306);
	nand gate_anoymous_9_n1154 (anoymous_9_n1154, anoymous_9_n932, anoymous_9_n931);
	or gate_anoymous_9_n930 (anoymous_9_n930, anoymous_9_n23, anoymous_9_n1306);
	or gate_anoymous_9_n929 (anoymous_9_n929, anoymous_9_n21, anoymous_9_n1305);
	nand gate_anoymous_9_n1153 (anoymous_9_n1153, anoymous_9_n930, anoymous_9_n929);
	or gate_anoymous_9_n928 (anoymous_9_n928, anoymous_9_n23, anoymous_9_n1305);
	or gate_anoymous_9_n927 (anoymous_9_n927, anoymous_9_n21, anoymous_9_n1304);
	nand gate_anoymous_9_n1152 (anoymous_9_n1152, anoymous_9_n928, anoymous_9_n927);
	or gate_anoymous_9_n926 (anoymous_9_n926, anoymous_9_n23, anoymous_9_n1304);
	or gate_anoymous_9_n925 (anoymous_9_n925, anoymous_9_n21, anoymous_9_n1303);
	nand gate_anoymous_9_n1151 (anoymous_9_n1151, anoymous_9_n926, anoymous_9_n925);
	or gate_anoymous_9_n924 (anoymous_9_n924, anoymous_9_n23, anoymous_9_n1303);
	or gate_anoymous_9_n923 (anoymous_9_n923, anoymous_9_n21, anoymous_9_n1302);
	nand gate_anoymous_9_n1150 (anoymous_9_n1150, anoymous_9_n924, anoymous_9_n923);
	or gate_anoymous_9_n922 (anoymous_9_n922, anoymous_9_n23, anoymous_9_n1302);
	or gate_anoymous_9_n921 (anoymous_9_n921, anoymous_9_n22, anoymous_9_n1301);
	nand gate_anoymous_9_n1149 (anoymous_9_n1149, anoymous_9_n922, anoymous_9_n921);
	or gate_anoymous_9_n920 (anoymous_9_n920, anoymous_9_n24, anoymous_9_n1301);
	or gate_anoymous_9_n919 (anoymous_9_n919, anoymous_9_n22, anoymous_9_n1300);
	nand gate_anoymous_9_n1148 (anoymous_9_n1148, anoymous_9_n920, anoymous_9_n919);
	or gate_anoymous_9_n918 (anoymous_9_n918, anoymous_9_n24, anoymous_9_n1300);
	or gate_anoymous_9_n917 (anoymous_9_n917, anoymous_9_n22, anoymous_9_n1299);
	nand gate_anoymous_9_n1147 (anoymous_9_n1147, anoymous_9_n918, anoymous_9_n917);
	or gate_anoymous_9_n916 (anoymous_9_n916, anoymous_9_n24, anoymous_9_n1299);
	or gate_anoymous_9_n915 (anoymous_9_n915, anoymous_9_n22, anoymous_9_n1298);
	nand gate_anoymous_9_n1146 (anoymous_9_n1146, anoymous_9_n916, anoymous_9_n915);
	or gate_anoymous_9_n914 (anoymous_9_n914, anoymous_9_n24, anoymous_9_n1298);
	or gate_anoymous_9_n913 (anoymous_9_n913, anoymous_9_n22, anoymous_9_n1297);
	nand gate_anoymous_9_n1145 (anoymous_9_n1145, anoymous_9_n914, anoymous_9_n913);
	or gate_anoymous_9_n912 (anoymous_9_n912, anoymous_9_n24, anoymous_9_n1297);
	or gate_anoymous_9_n911 (anoymous_9_n911, anoymous_9_n22, anoymous_9_n1296);
	nand gate_anoymous_9_n1144 (anoymous_9_n1144, anoymous_9_n912, anoymous_9_n911);
	or gate_anoymous_9_n910 (anoymous_9_n910, anoymous_9_n24, anoymous_9_n1296);
	or gate_anoymous_9_n909 (anoymous_9_n909, anoymous_9_n22, anoymous_9_n1295);
	nand gate_anoymous_9_n1143 (anoymous_9_n1143, anoymous_9_n910, anoymous_9_n909);
	or gate_anoymous_9_n908 (anoymous_9_n908, anoymous_9_n24, anoymous_9_n1295);
	or gate_anoymous_9_n907 (anoymous_9_n907, anoymous_9_n22, anoymous_9_n1408);
	nand gate_anoymous_9_n1142 (anoymous_9_n1142, anoymous_9_n908, anoymous_9_n907);
	and gate_anoymous_9_n906 (anoymous_9_n906, anoymous_9_n24, anoymous_9_n22);
	or gate_anoymous_9_n1141 (anoymous_9_n1141, anoymous_9_n1408, anoymous_9_n906);
	or gate_anoymous_9_n905 (anoymous_9_n905, anoymous_9_n22, anoymous_9_n1311);
	or gate_anoymous_9_n904 (anoymous_9_n904, anoymous_9_n24, anoymous_9_n1408);
	nand gate_anoymous_9_n1056 (anoymous_9_n1056, anoymous_9_n905, anoymous_9_n904);
	or gate_anoymous_9_n1294 (anoymous_9_n1294, anoymous_9_n49, anoymous_9_n1407);
	xnor gate_anoymous_9_n1293 (anoymous_9_n1293, anoymous_9_n49, anoymous_9_n25);
	xnor gate_anoymous_9_n1292 (anoymous_9_n1292, anoymous_9_n1377, anoymous_9_n25);
	xnor gate_anoymous_9_n1291 (anoymous_9_n1291, anoymous_9_n1376, anoymous_9_n25);
	xnor gate_anoymous_9_n1290 (anoymous_9_n1290, anoymous_9_n1375, anoymous_9_n25);
	xnor gate_anoymous_9_n1289 (anoymous_9_n1289, anoymous_9_n1374, anoymous_9_n25);
	xnor gate_anoymous_9_n1288 (anoymous_9_n1288, anoymous_9_n1373, anoymous_9_n25);
	xnor gate_anoymous_9_n1287 (anoymous_9_n1287, anoymous_9_n1372, anoymous_9_n25);
	xnor gate_anoymous_9_n1286 (anoymous_9_n1286, anoymous_9_n1371, anoymous_9_n25);
	xnor gate_anoymous_9_n1285 (anoymous_9_n1285, anoymous_9_n1370, anoymous_9_n25);
	xnor gate_anoymous_9_n1284 (anoymous_9_n1284, anoymous_9_n1369, anoymous_9_n25);
	xnor gate_anoymous_9_n1283 (anoymous_9_n1283, anoymous_9_n1368, anoymous_9_n25);
	xnor gate_anoymous_9_n1282 (anoymous_9_n1282, anoymous_9_n1367, anoymous_9_n25);
	xnor gate_anoymous_9_n1281 (anoymous_9_n1281, anoymous_9_n1366, anoymous_9_n25);
	xnor gate_anoymous_9_n1280 (anoymous_9_n1280, anoymous_9_n1365, anoymous_9_n25);
	xnor gate_anoymous_9_n1279 (anoymous_9_n1279, anoymous_9_n1364, anoymous_9_n25);
	xnor gate_anoymous_9_n1278 (anoymous_9_n1278, anoymous_9_n1363, anoymous_9_n25);
	not gate_anoymous_9_n902 (anoymous_9_n902, anoymous_9_n27);
	and gate_anoymous_9_n1140 (anoymous_9_n1140, anoymous_9_n49, anoymous_9_n902);
	or gate_anoymous_9_n901 (anoymous_9_n901, anoymous_9_n29, anoymous_9_n1293);
	or gate_anoymous_9_n900 (anoymous_9_n900, anoymous_9_n27, anoymous_9_n1292);
	nand gate_anoymous_9_n1139 (anoymous_9_n1139, anoymous_9_n901, anoymous_9_n900);
	or gate_anoymous_9_n899 (anoymous_9_n899, anoymous_9_n29, anoymous_9_n1292);
	or gate_anoymous_9_n898 (anoymous_9_n898, anoymous_9_n27, anoymous_9_n1291);
	nand gate_anoymous_9_n1138 (anoymous_9_n1138, anoymous_9_n899, anoymous_9_n898);
	or gate_anoymous_9_n897 (anoymous_9_n897, anoymous_9_n29, anoymous_9_n1291);
	or gate_anoymous_9_n896 (anoymous_9_n896, anoymous_9_n27, anoymous_9_n1290);
	nand gate_anoymous_9_n1137 (anoymous_9_n1137, anoymous_9_n897, anoymous_9_n896);
	or gate_anoymous_9_n895 (anoymous_9_n895, anoymous_9_n29, anoymous_9_n1290);
	or gate_anoymous_9_n894 (anoymous_9_n894, anoymous_9_n27, anoymous_9_n1289);
	nand gate_anoymous_9_n1136 (anoymous_9_n1136, anoymous_9_n895, anoymous_9_n894);
	or gate_anoymous_9_n893 (anoymous_9_n893, anoymous_9_n29, anoymous_9_n1289);
	or gate_anoymous_9_n892 (anoymous_9_n892, anoymous_9_n27, anoymous_9_n1288);
	nand gate_anoymous_9_n1135 (anoymous_9_n1135, anoymous_9_n893, anoymous_9_n892);
	or gate_anoymous_9_n891 (anoymous_9_n891, anoymous_9_n29, anoymous_9_n1288);
	or gate_anoymous_9_n890 (anoymous_9_n890, anoymous_9_n27, anoymous_9_n1287);
	nand gate_anoymous_9_n1134 (anoymous_9_n1134, anoymous_9_n891, anoymous_9_n890);
	or gate_anoymous_9_n889 (anoymous_9_n889, anoymous_9_n29, anoymous_9_n1287);
	or gate_anoymous_9_n888 (anoymous_9_n888, anoymous_9_n27, anoymous_9_n1286);
	nand gate_anoymous_9_n1133 (anoymous_9_n1133, anoymous_9_n889, anoymous_9_n888);
	or gate_anoymous_9_n887 (anoymous_9_n887, anoymous_9_n29, anoymous_9_n1286);
	or gate_anoymous_9_n886 (anoymous_9_n886, anoymous_9_n27, anoymous_9_n1285);
	nand gate_anoymous_9_n1132 (anoymous_9_n1132, anoymous_9_n887, anoymous_9_n886);
	or gate_anoymous_9_n885 (anoymous_9_n885, anoymous_9_n29, anoymous_9_n1285);
	or gate_anoymous_9_n884 (anoymous_9_n884, anoymous_9_n28, anoymous_9_n1284);
	nand gate_anoymous_9_n1131 (anoymous_9_n1131, anoymous_9_n885, anoymous_9_n884);
	or gate_anoymous_9_n883 (anoymous_9_n883, anoymous_9_n30, anoymous_9_n1284);
	or gate_anoymous_9_n882 (anoymous_9_n882, anoymous_9_n28, anoymous_9_n1283);
	nand gate_anoymous_9_n1130 (anoymous_9_n1130, anoymous_9_n883, anoymous_9_n882);
	or gate_anoymous_9_n881 (anoymous_9_n881, anoymous_9_n30, anoymous_9_n1283);
	or gate_anoymous_9_n880 (anoymous_9_n880, anoymous_9_n28, anoymous_9_n1282);
	nand gate_anoymous_9_n1129 (anoymous_9_n1129, anoymous_9_n881, anoymous_9_n880);
	or gate_anoymous_9_n879 (anoymous_9_n879, anoymous_9_n30, anoymous_9_n1282);
	or gate_anoymous_9_n878 (anoymous_9_n878, anoymous_9_n28, anoymous_9_n1281);
	nand gate_anoymous_9_n1128 (anoymous_9_n1128, anoymous_9_n879, anoymous_9_n878);
	or gate_anoymous_9_n877 (anoymous_9_n877, anoymous_9_n30, anoymous_9_n1281);
	or gate_anoymous_9_n876 (anoymous_9_n876, anoymous_9_n28, anoymous_9_n1280);
	nand gate_anoymous_9_n1127 (anoymous_9_n1127, anoymous_9_n877, anoymous_9_n876);
	or gate_anoymous_9_n875 (anoymous_9_n875, anoymous_9_n30, anoymous_9_n1280);
	or gate_anoymous_9_n874 (anoymous_9_n874, anoymous_9_n28, anoymous_9_n1279);
	nand gate_anoymous_9_n1126 (anoymous_9_n1126, anoymous_9_n875, anoymous_9_n874);
	or gate_anoymous_9_n873 (anoymous_9_n873, anoymous_9_n30, anoymous_9_n1279);
	or gate_anoymous_9_n872 (anoymous_9_n872, anoymous_9_n28, anoymous_9_n1278);
	nand gate_anoymous_9_n1125 (anoymous_9_n1125, anoymous_9_n873, anoymous_9_n872);
	or gate_anoymous_9_n871 (anoymous_9_n871, anoymous_9_n30, anoymous_9_n1278);
	or gate_anoymous_9_n870 (anoymous_9_n870, anoymous_9_n28, anoymous_9_n1407);
	nand gate_anoymous_9_n1124 (anoymous_9_n1124, anoymous_9_n871, anoymous_9_n870);
	and gate_anoymous_9_n869 (anoymous_9_n869, anoymous_9_n30, anoymous_9_n28);
	or gate_anoymous_9_n1123 (anoymous_9_n1123, anoymous_9_n1407, anoymous_9_n869);
	or gate_anoymous_9_n868 (anoymous_9_n868, anoymous_9_n28, anoymous_9_n1294);
	or gate_anoymous_9_n867 (anoymous_9_n867, anoymous_9_n30, anoymous_9_n1407);
	nand gate_anoymous_9_n1055 (anoymous_9_n1055, anoymous_9_n868, anoymous_9_n867);
	or gate_anoymous_9_n1277 (anoymous_9_n1277, anoymous_9_n49, anoymous_9_n1406);
	xnor gate_anoymous_9_n1276 (anoymous_9_n1276, anoymous_9_n49, anoymous_9_n31);
	xnor gate_anoymous_9_n1275 (anoymous_9_n1275, anoymous_9_n1377, anoymous_9_n31);
	xnor gate_anoymous_9_n1274 (anoymous_9_n1274, anoymous_9_n1376, anoymous_9_n31);
	xnor gate_anoymous_9_n1273 (anoymous_9_n1273, anoymous_9_n1375, anoymous_9_n31);
	xnor gate_anoymous_9_n1272 (anoymous_9_n1272, anoymous_9_n1374, anoymous_9_n31);
	xnor gate_anoymous_9_n1271 (anoymous_9_n1271, anoymous_9_n1373, anoymous_9_n31);
	xnor gate_anoymous_9_n1270 (anoymous_9_n1270, anoymous_9_n1372, anoymous_9_n31);
	xnor gate_anoymous_9_n1269 (anoymous_9_n1269, anoymous_9_n1371, anoymous_9_n31);
	xnor gate_anoymous_9_n1268 (anoymous_9_n1268, anoymous_9_n1370, anoymous_9_n31);
	xnor gate_anoymous_9_n1267 (anoymous_9_n1267, anoymous_9_n1369, anoymous_9_n31);
	xnor gate_anoymous_9_n1266 (anoymous_9_n1266, anoymous_9_n1368, anoymous_9_n31);
	xnor gate_anoymous_9_n1265 (anoymous_9_n1265, anoymous_9_n1367, anoymous_9_n31);
	xnor gate_anoymous_9_n1264 (anoymous_9_n1264, anoymous_9_n1366, anoymous_9_n31);
	xnor gate_anoymous_9_n1263 (anoymous_9_n1263, anoymous_9_n1365, anoymous_9_n31);
	xnor gate_anoymous_9_n1262 (anoymous_9_n1262, anoymous_9_n1364, anoymous_9_n31);
	xnor gate_anoymous_9_n1261 (anoymous_9_n1261, anoymous_9_n1363, anoymous_9_n31);
	not gate_anoymous_9_n865 (anoymous_9_n865, anoymous_9_n33);
	and gate_anoymous_9_n1122 (anoymous_9_n1122, anoymous_9_n49, anoymous_9_n865);
	or gate_anoymous_9_n864 (anoymous_9_n864, anoymous_9_n35, anoymous_9_n1276);
	or gate_anoymous_9_n863 (anoymous_9_n863, anoymous_9_n33, anoymous_9_n1275);
	nand gate_anoymous_9_n1121 (anoymous_9_n1121, anoymous_9_n864, anoymous_9_n863);
	or gate_anoymous_9_n862 (anoymous_9_n862, anoymous_9_n35, anoymous_9_n1275);
	or gate_anoymous_9_n861 (anoymous_9_n861, anoymous_9_n33, anoymous_9_n1274);
	nand gate_anoymous_9_n1120 (anoymous_9_n1120, anoymous_9_n862, anoymous_9_n861);
	or gate_anoymous_9_n860 (anoymous_9_n860, anoymous_9_n35, anoymous_9_n1274);
	or gate_anoymous_9_n859 (anoymous_9_n859, anoymous_9_n33, anoymous_9_n1273);
	nand gate_anoymous_9_n1119 (anoymous_9_n1119, anoymous_9_n860, anoymous_9_n859);
	or gate_anoymous_9_n858 (anoymous_9_n858, anoymous_9_n35, anoymous_9_n1273);
	or gate_anoymous_9_n857 (anoymous_9_n857, anoymous_9_n33, anoymous_9_n1272);
	nand gate_anoymous_9_n1118 (anoymous_9_n1118, anoymous_9_n858, anoymous_9_n857);
	or gate_anoymous_9_n856 (anoymous_9_n856, anoymous_9_n35, anoymous_9_n1272);
	or gate_anoymous_9_n855 (anoymous_9_n855, anoymous_9_n33, anoymous_9_n1271);
	nand gate_anoymous_9_n1117 (anoymous_9_n1117, anoymous_9_n856, anoymous_9_n855);
	or gate_anoymous_9_n854 (anoymous_9_n854, anoymous_9_n35, anoymous_9_n1271);
	or gate_anoymous_9_n853 (anoymous_9_n853, anoymous_9_n33, anoymous_9_n1270);
	nand gate_anoymous_9_n1116 (anoymous_9_n1116, anoymous_9_n854, anoymous_9_n853);
	or gate_anoymous_9_n852 (anoymous_9_n852, anoymous_9_n35, anoymous_9_n1270);
	or gate_anoymous_9_n851 (anoymous_9_n851, anoymous_9_n33, anoymous_9_n1269);
	nand gate_anoymous_9_n1115 (anoymous_9_n1115, anoymous_9_n852, anoymous_9_n851);
	or gate_anoymous_9_n850 (anoymous_9_n850, anoymous_9_n35, anoymous_9_n1269);
	or gate_anoymous_9_n849 (anoymous_9_n849, anoymous_9_n33, anoymous_9_n1268);
	nand gate_anoymous_9_n1114 (anoymous_9_n1114, anoymous_9_n850, anoymous_9_n849);
	or gate_anoymous_9_n848 (anoymous_9_n848, anoymous_9_n35, anoymous_9_n1268);
	or gate_anoymous_9_n847 (anoymous_9_n847, anoymous_9_n34, anoymous_9_n1267);
	nand gate_anoymous_9_n1113 (anoymous_9_n1113, anoymous_9_n848, anoymous_9_n847);
	or gate_anoymous_9_n846 (anoymous_9_n846, anoymous_9_n36, anoymous_9_n1267);
	or gate_anoymous_9_n845 (anoymous_9_n845, anoymous_9_n34, anoymous_9_n1266);
	nand gate_anoymous_9_n1112 (anoymous_9_n1112, anoymous_9_n846, anoymous_9_n845);
	or gate_anoymous_9_n844 (anoymous_9_n844, anoymous_9_n36, anoymous_9_n1266);
	or gate_anoymous_9_n843 (anoymous_9_n843, anoymous_9_n34, anoymous_9_n1265);
	nand gate_anoymous_9_n1111 (anoymous_9_n1111, anoymous_9_n844, anoymous_9_n843);
	or gate_anoymous_9_n842 (anoymous_9_n842, anoymous_9_n36, anoymous_9_n1265);
	or gate_anoymous_9_n841 (anoymous_9_n841, anoymous_9_n34, anoymous_9_n1264);
	nand gate_anoymous_9_n1110 (anoymous_9_n1110, anoymous_9_n842, anoymous_9_n841);
	or gate_anoymous_9_n840 (anoymous_9_n840, anoymous_9_n36, anoymous_9_n1264);
	or gate_anoymous_9_n839 (anoymous_9_n839, anoymous_9_n34, anoymous_9_n1263);
	nand gate_anoymous_9_n1109 (anoymous_9_n1109, anoymous_9_n840, anoymous_9_n839);
	or gate_anoymous_9_n838 (anoymous_9_n838, anoymous_9_n36, anoymous_9_n1263);
	or gate_anoymous_9_n837 (anoymous_9_n837, anoymous_9_n34, anoymous_9_n1262);
	nand gate_anoymous_9_n1108 (anoymous_9_n1108, anoymous_9_n838, anoymous_9_n837);
	or gate_anoymous_9_n836 (anoymous_9_n836, anoymous_9_n36, anoymous_9_n1262);
	or gate_anoymous_9_n835 (anoymous_9_n835, anoymous_9_n34, anoymous_9_n1261);
	nand gate_anoymous_9_n1107 (anoymous_9_n1107, anoymous_9_n836, anoymous_9_n835);
	or gate_anoymous_9_n834 (anoymous_9_n834, anoymous_9_n36, anoymous_9_n1261);
	or gate_anoymous_9_n833 (anoymous_9_n833, anoymous_9_n34, anoymous_9_n1406);
	nand gate_anoymous_9_n1106 (anoymous_9_n1106, anoymous_9_n834, anoymous_9_n833);
	and gate_anoymous_9_n832 (anoymous_9_n832, anoymous_9_n36, anoymous_9_n34);
	or gate_anoymous_9_n1105 (anoymous_9_n1105, anoymous_9_n1406, anoymous_9_n832);
	or gate_anoymous_9_n831 (anoymous_9_n831, anoymous_9_n34, anoymous_9_n1277);
	or gate_anoymous_9_n830 (anoymous_9_n830, anoymous_9_n36, anoymous_9_n1406);
	nand gate_anoymous_9_n1054 (anoymous_9_n1054, anoymous_9_n831, anoymous_9_n830);
	or gate_anoymous_9_n1260 (anoymous_9_n1260, anoymous_9_n49, anoymous_9_n1405);
	xnor gate_anoymous_9_n1259 (anoymous_9_n1259, anoymous_9_n49, anoymous_9_n37);
	xnor gate_anoymous_9_n1258 (anoymous_9_n1258, anoymous_9_n1377, anoymous_9_n37);
	xnor gate_anoymous_9_n1257 (anoymous_9_n1257, anoymous_9_n1376, anoymous_9_n37);
	xnor gate_anoymous_9_n1256 (anoymous_9_n1256, anoymous_9_n1375, anoymous_9_n37);
	xnor gate_anoymous_9_n1255 (anoymous_9_n1255, anoymous_9_n1374, anoymous_9_n37);
	xnor gate_anoymous_9_n1254 (anoymous_9_n1254, anoymous_9_n1373, anoymous_9_n37);
	xnor gate_anoymous_9_n1253 (anoymous_9_n1253, anoymous_9_n1372, anoymous_9_n37);
	xnor gate_anoymous_9_n1252 (anoymous_9_n1252, anoymous_9_n1371, anoymous_9_n37);
	xnor gate_anoymous_9_n1251 (anoymous_9_n1251, anoymous_9_n1370, anoymous_9_n37);
	xnor gate_anoymous_9_n1250 (anoymous_9_n1250, anoymous_9_n1369, anoymous_9_n37);
	xnor gate_anoymous_9_n1249 (anoymous_9_n1249, anoymous_9_n1368, anoymous_9_n37);
	xnor gate_anoymous_9_n1248 (anoymous_9_n1248, anoymous_9_n1367, anoymous_9_n37);
	xnor gate_anoymous_9_n1247 (anoymous_9_n1247, anoymous_9_n1366, anoymous_9_n37);
	xnor gate_anoymous_9_n1246 (anoymous_9_n1246, anoymous_9_n1365, anoymous_9_n37);
	xnor gate_anoymous_9_n1245 (anoymous_9_n1245, anoymous_9_n1364, anoymous_9_n37);
	xnor gate_anoymous_9_n1244 (anoymous_9_n1244, anoymous_9_n1363, anoymous_9_n37);
	not gate_anoymous_9_n828 (anoymous_9_n828, anoymous_9_n39);
	and gate_anoymous_9_n1104 (anoymous_9_n1104, anoymous_9_n49, anoymous_9_n828);
	or gate_anoymous_9_n827 (anoymous_9_n827, anoymous_9_n41, anoymous_9_n1259);
	or gate_anoymous_9_n826 (anoymous_9_n826, anoymous_9_n39, anoymous_9_n1258);
	nand gate_anoymous_9_n1103 (anoymous_9_n1103, anoymous_9_n827, anoymous_9_n826);
	or gate_anoymous_9_n825 (anoymous_9_n825, anoymous_9_n41, anoymous_9_n1258);
	or gate_anoymous_9_n824 (anoymous_9_n824, anoymous_9_n39, anoymous_9_n1257);
	nand gate_anoymous_9_n1102 (anoymous_9_n1102, anoymous_9_n825, anoymous_9_n824);
	or gate_anoymous_9_n823 (anoymous_9_n823, anoymous_9_n41, anoymous_9_n1257);
	or gate_anoymous_9_n822 (anoymous_9_n822, anoymous_9_n39, anoymous_9_n1256);
	nand gate_anoymous_9_n1101 (anoymous_9_n1101, anoymous_9_n823, anoymous_9_n822);
	or gate_anoymous_9_n821 (anoymous_9_n821, anoymous_9_n41, anoymous_9_n1256);
	or gate_anoymous_9_n820 (anoymous_9_n820, anoymous_9_n39, anoymous_9_n1255);
	nand gate_anoymous_9_n1100 (anoymous_9_n1100, anoymous_9_n821, anoymous_9_n820);
	or gate_anoymous_9_n819 (anoymous_9_n819, anoymous_9_n41, anoymous_9_n1255);
	or gate_anoymous_9_n818 (anoymous_9_n818, anoymous_9_n39, anoymous_9_n1254);
	nand gate_anoymous_9_n1099 (anoymous_9_n1099, anoymous_9_n819, anoymous_9_n818);
	or gate_anoymous_9_n817 (anoymous_9_n817, anoymous_9_n41, anoymous_9_n1254);
	or gate_anoymous_9_n816 (anoymous_9_n816, anoymous_9_n39, anoymous_9_n1253);
	nand gate_anoymous_9_n1098 (anoymous_9_n1098, anoymous_9_n817, anoymous_9_n816);
	or gate_anoymous_9_n815 (anoymous_9_n815, anoymous_9_n41, anoymous_9_n1253);
	or gate_anoymous_9_n814 (anoymous_9_n814, anoymous_9_n39, anoymous_9_n1252);
	nand gate_anoymous_9_n1097 (anoymous_9_n1097, anoymous_9_n815, anoymous_9_n814);
	or gate_anoymous_9_n813 (anoymous_9_n813, anoymous_9_n41, anoymous_9_n1252);
	or gate_anoymous_9_n812 (anoymous_9_n812, anoymous_9_n39, anoymous_9_n1251);
	nand gate_anoymous_9_n1096 (anoymous_9_n1096, anoymous_9_n813, anoymous_9_n812);
	or gate_anoymous_9_n811 (anoymous_9_n811, anoymous_9_n41, anoymous_9_n1251);
	or gate_anoymous_9_n810 (anoymous_9_n810, anoymous_9_n40, anoymous_9_n1250);
	nand gate_anoymous_9_n1095 (anoymous_9_n1095, anoymous_9_n811, anoymous_9_n810);
	or gate_anoymous_9_n809 (anoymous_9_n809, anoymous_9_n42, anoymous_9_n1250);
	or gate_anoymous_9_n808 (anoymous_9_n808, anoymous_9_n40, anoymous_9_n1249);
	nand gate_anoymous_9_n1094 (anoymous_9_n1094, anoymous_9_n809, anoymous_9_n808);
	or gate_anoymous_9_n807 (anoymous_9_n807, anoymous_9_n42, anoymous_9_n1249);
	or gate_anoymous_9_n806 (anoymous_9_n806, anoymous_9_n40, anoymous_9_n1248);
	nand gate_anoymous_9_n1093 (anoymous_9_n1093, anoymous_9_n807, anoymous_9_n806);
	or gate_anoymous_9_n805 (anoymous_9_n805, anoymous_9_n42, anoymous_9_n1248);
	or gate_anoymous_9_n804 (anoymous_9_n804, anoymous_9_n40, anoymous_9_n1247);
	nand gate_anoymous_9_n1092 (anoymous_9_n1092, anoymous_9_n805, anoymous_9_n804);
	or gate_anoymous_9_n803 (anoymous_9_n803, anoymous_9_n42, anoymous_9_n1247);
	or gate_anoymous_9_n802 (anoymous_9_n802, anoymous_9_n40, anoymous_9_n1246);
	nand gate_anoymous_9_n1091 (anoymous_9_n1091, anoymous_9_n803, anoymous_9_n802);
	or gate_anoymous_9_n801 (anoymous_9_n801, anoymous_9_n42, anoymous_9_n1246);
	or gate_anoymous_9_n800 (anoymous_9_n800, anoymous_9_n40, anoymous_9_n1245);
	nand gate_anoymous_9_n1090 (anoymous_9_n1090, anoymous_9_n801, anoymous_9_n800);
	or gate_anoymous_9_n799 (anoymous_9_n799, anoymous_9_n42, anoymous_9_n1245);
	or gate_anoymous_9_n798 (anoymous_9_n798, anoymous_9_n40, anoymous_9_n1244);
	nand gate_anoymous_9_n1089 (anoymous_9_n1089, anoymous_9_n799, anoymous_9_n798);
	or gate_anoymous_9_n797 (anoymous_9_n797, anoymous_9_n42, anoymous_9_n1244);
	or gate_anoymous_9_n796 (anoymous_9_n796, anoymous_9_n40, anoymous_9_n1405);
	nand gate_anoymous_9_n1088 (anoymous_9_n1088, anoymous_9_n797, anoymous_9_n796);
	and gate_anoymous_9_n795 (anoymous_9_n795, anoymous_9_n42, anoymous_9_n40);
	or gate_anoymous_9_n1087 (anoymous_9_n1087, anoymous_9_n1405, anoymous_9_n795);
	or gate_anoymous_9_n794 (anoymous_9_n794, anoymous_9_n40, anoymous_9_n1260);
	or gate_anoymous_9_n793 (anoymous_9_n793, anoymous_9_n42, anoymous_9_n1405);
	nand gate_anoymous_9_n1053 (anoymous_9_n1053, anoymous_9_n794, anoymous_9_n793);
	or gate_anoymous_9_n1243 (anoymous_9_n1243, anoymous_9_n49, anoymous_9_n1404);
	xnor gate_anoymous_9_n1242 (anoymous_9_n1242, anoymous_9_n49, anoymous_9_n43);
	xnor gate_anoymous_9_n1241 (anoymous_9_n1241, anoymous_9_n1377, anoymous_9_n43);
	xnor gate_anoymous_9_n1240 (anoymous_9_n1240, anoymous_9_n1376, anoymous_9_n43);
	xnor gate_anoymous_9_n1239 (anoymous_9_n1239, anoymous_9_n1375, anoymous_9_n43);
	xnor gate_anoymous_9_n1238 (anoymous_9_n1238, anoymous_9_n1374, anoymous_9_n43);
	xnor gate_anoymous_9_n1237 (anoymous_9_n1237, anoymous_9_n1373, anoymous_9_n43);
	xnor gate_anoymous_9_n1236 (anoymous_9_n1236, anoymous_9_n1372, anoymous_9_n43);
	xnor gate_anoymous_9_n1235 (anoymous_9_n1235, anoymous_9_n1371, anoymous_9_n43);
	xnor gate_anoymous_9_n1234 (anoymous_9_n1234, anoymous_9_n1370, anoymous_9_n43);
	xnor gate_anoymous_9_n1233 (anoymous_9_n1233, anoymous_9_n1369, anoymous_9_n43);
	xnor gate_anoymous_9_n1232 (anoymous_9_n1232, anoymous_9_n1368, anoymous_9_n43);
	xnor gate_anoymous_9_n1231 (anoymous_9_n1231, anoymous_9_n1367, anoymous_9_n43);
	xnor gate_anoymous_9_n1230 (anoymous_9_n1230, anoymous_9_n1366, anoymous_9_n43);
	xnor gate_anoymous_9_n1229 (anoymous_9_n1229, anoymous_9_n1365, anoymous_9_n43);
	xnor gate_anoymous_9_n1228 (anoymous_9_n1228, anoymous_9_n1364, anoymous_9_n43);
	xnor gate_anoymous_9_n1227 (anoymous_9_n1227, anoymous_9_n1363, anoymous_9_n43);
	not gate_anoymous_9_n791 (anoymous_9_n791, anoymous_9_n45);
	and gate_anoymous_9_n1086 (anoymous_9_n1086, anoymous_9_n49, anoymous_9_n791);
	or gate_anoymous_9_n790 (anoymous_9_n790, anoymous_9_n47, anoymous_9_n1242);
	or gate_anoymous_9_n789 (anoymous_9_n789, anoymous_9_n45, anoymous_9_n1241);
	nand gate_anoymous_9_n1085 (anoymous_9_n1085, anoymous_9_n790, anoymous_9_n789);
	or gate_anoymous_9_n788 (anoymous_9_n788, anoymous_9_n47, anoymous_9_n1241);
	or gate_anoymous_9_n787 (anoymous_9_n787, anoymous_9_n45, anoymous_9_n1240);
	nand gate_anoymous_9_n1084 (anoymous_9_n1084, anoymous_9_n788, anoymous_9_n787);
	or gate_anoymous_9_n786 (anoymous_9_n786, anoymous_9_n47, anoymous_9_n1240);
	or gate_anoymous_9_n785 (anoymous_9_n785, anoymous_9_n45, anoymous_9_n1239);
	nand gate_anoymous_9_n1083 (anoymous_9_n1083, anoymous_9_n786, anoymous_9_n785);
	or gate_anoymous_9_n784 (anoymous_9_n784, anoymous_9_n47, anoymous_9_n1239);
	or gate_anoymous_9_n783 (anoymous_9_n783, anoymous_9_n45, anoymous_9_n1238);
	nand gate_anoymous_9_n1082 (anoymous_9_n1082, anoymous_9_n784, anoymous_9_n783);
	or gate_anoymous_9_n782 (anoymous_9_n782, anoymous_9_n47, anoymous_9_n1238);
	or gate_anoymous_9_n781 (anoymous_9_n781, anoymous_9_n45, anoymous_9_n1237);
	nand gate_anoymous_9_n1081 (anoymous_9_n1081, anoymous_9_n782, anoymous_9_n781);
	or gate_anoymous_9_n780 (anoymous_9_n780, anoymous_9_n47, anoymous_9_n1237);
	or gate_anoymous_9_n779 (anoymous_9_n779, anoymous_9_n45, anoymous_9_n1236);
	nand gate_anoymous_9_n1080 (anoymous_9_n1080, anoymous_9_n780, anoymous_9_n779);
	or gate_anoymous_9_n778 (anoymous_9_n778, anoymous_9_n47, anoymous_9_n1236);
	or gate_anoymous_9_n777 (anoymous_9_n777, anoymous_9_n45, anoymous_9_n1235);
	nand gate_anoymous_9_n1079 (anoymous_9_n1079, anoymous_9_n778, anoymous_9_n777);
	or gate_anoymous_9_n776 (anoymous_9_n776, anoymous_9_n47, anoymous_9_n1235);
	or gate_anoymous_9_n775 (anoymous_9_n775, anoymous_9_n45, anoymous_9_n1234);
	nand gate_anoymous_9_n1078 (anoymous_9_n1078, anoymous_9_n776, anoymous_9_n775);
	or gate_anoymous_9_n774 (anoymous_9_n774, anoymous_9_n47, anoymous_9_n1234);
	or gate_anoymous_9_n773 (anoymous_9_n773, anoymous_9_n46, anoymous_9_n1233);
	nand gate_anoymous_9_n1077 (anoymous_9_n1077, anoymous_9_n774, anoymous_9_n773);
	or gate_anoymous_9_n772 (anoymous_9_n772, anoymous_9_n48, anoymous_9_n1233);
	or gate_anoymous_9_n771 (anoymous_9_n771, anoymous_9_n46, anoymous_9_n1232);
	nand gate_anoymous_9_n1076 (anoymous_9_n1076, anoymous_9_n772, anoymous_9_n771);
	or gate_anoymous_9_n770 (anoymous_9_n770, anoymous_9_n48, anoymous_9_n1232);
	or gate_anoymous_9_n769 (anoymous_9_n769, anoymous_9_n46, anoymous_9_n1231);
	nand gate_anoymous_9_n1075 (anoymous_9_n1075, anoymous_9_n770, anoymous_9_n769);
	or gate_anoymous_9_n768 (anoymous_9_n768, anoymous_9_n48, anoymous_9_n1231);
	or gate_anoymous_9_n767 (anoymous_9_n767, anoymous_9_n46, anoymous_9_n1230);
	nand gate_anoymous_9_n1074 (anoymous_9_n1074, anoymous_9_n768, anoymous_9_n767);
	or gate_anoymous_9_n766 (anoymous_9_n766, anoymous_9_n48, anoymous_9_n1230);
	or gate_anoymous_9_n765 (anoymous_9_n765, anoymous_9_n46, anoymous_9_n1229);
	nand gate_anoymous_9_n1073 (anoymous_9_n1073, anoymous_9_n766, anoymous_9_n765);
	or gate_anoymous_9_n764 (anoymous_9_n764, anoymous_9_n48, anoymous_9_n1229);
	or gate_anoymous_9_n763 (anoymous_9_n763, anoymous_9_n46, anoymous_9_n1228);
	nand gate_anoymous_9_n1072 (anoymous_9_n1072, anoymous_9_n764, anoymous_9_n763);
	or gate_anoymous_9_n762 (anoymous_9_n762, anoymous_9_n48, anoymous_9_n1228);
	or gate_anoymous_9_n761 (anoymous_9_n761, anoymous_9_n46, anoymous_9_n1227);
	nand gate_anoymous_9_n1071 (anoymous_9_n1071, anoymous_9_n762, anoymous_9_n761);
	or gate_anoymous_9_n760 (anoymous_9_n760, anoymous_9_n48, anoymous_9_n1227);
	or gate_anoymous_9_n759 (anoymous_9_n759, anoymous_9_n46, anoymous_9_n1404);
	nand gate_anoymous_9_n1070 (anoymous_9_n1070, anoymous_9_n760, anoymous_9_n759);
	and gate_anoymous_9_n758 (anoymous_9_n758, anoymous_9_n48, anoymous_9_n46);
	or gate_anoymous_9_n1069 (anoymous_9_n1069, anoymous_9_n1404, anoymous_9_n758);
	or gate_anoymous_9_n757 (anoymous_9_n757, anoymous_9_n46, anoymous_9_n1243);
	or gate_anoymous_9_n756 (anoymous_9_n756, anoymous_9_n48, anoymous_9_n1404);
	nand gate_anoymous_9_n1052 (anoymous_9_n1052, anoymous_9_n757, anoymous_9_n756);
	not gate_anoymous_9_n1226 (anoymous_9_n1226, anoymous_9_n1377);
	not gate_anoymous_9_n1225 (anoymous_9_n1225, anoymous_9_n1376);
	not gate_anoymous_9_n1224 (anoymous_9_n1224, anoymous_9_n1375);
	not gate_anoymous_9_n1223 (anoymous_9_n1223, anoymous_9_n1374);
	not gate_anoymous_9_n1222 (anoymous_9_n1222, anoymous_9_n1373);
	not gate_anoymous_9_n1221 (anoymous_9_n1221, anoymous_9_n1372);
	not gate_anoymous_9_n1220 (anoymous_9_n1220, anoymous_9_n1371);
	not gate_anoymous_9_n1219 (anoymous_9_n1219, anoymous_9_n1370);
	not gate_anoymous_9_n1218 (anoymous_9_n1218, anoymous_9_n1369);
	not gate_anoymous_9_n1217 (anoymous_9_n1217, anoymous_9_n1368);
	not gate_anoymous_9_n1216 (anoymous_9_n1216, anoymous_9_n1367);
	not gate_anoymous_9_n1215 (anoymous_9_n1215, anoymous_9_n1366);
	not gate_anoymous_9_n1214 (anoymous_9_n1214, anoymous_9_n1365);
	not gate_anoymous_9_n1213 (anoymous_9_n1213, anoymous_9_n1364);
	not gate_anoymous_9_n1212 (anoymous_9_n1212, anoymous_9_n1363);
	not gate_anoymous_9_n755 (anoymous_9_n755, anoymous_9_n1395);
	and gate_anoymous_9_n1068 (anoymous_9_n1068, anoymous_9_n49, anoymous_9_n755);
	nor gate_anoymous_9_n458 (anoymous_9_n458, anoymous_9_n1226, anoymous_9_n1395);
	nor gate_anoymous_9_n1067 (anoymous_9_n1067, anoymous_9_n1225, anoymous_9_n1395);
	nor gate_anoymous_9_n1066 (anoymous_9_n1066, anoymous_9_n1224, anoymous_9_n1395);
	nor gate_anoymous_9_n386 (anoymous_9_n386, anoymous_9_n1223, anoymous_9_n1395);
	nor gate_anoymous_9_n1065 (anoymous_9_n1065, anoymous_9_n1222, anoymous_9_n1395);
	nor gate_anoymous_9_n324 (anoymous_9_n324, anoymous_9_n1221, anoymous_9_n1395);
	nor gate_anoymous_9_n1064 (anoymous_9_n1064, anoymous_9_n1220, anoymous_9_n1395);
	nor gate_anoymous_9_n272 (anoymous_9_n272, anoymous_9_n1219, anoymous_9_n1395);
	nor gate_anoymous_9_n1063 (anoymous_9_n1063, anoymous_9_n1218, anoymous_9_n1395);
	nor gate_anoymous_9_n230 (anoymous_9_n230, anoymous_9_n1217, anoymous_9_n1395);
	nor gate_anoymous_9_n1062 (anoymous_9_n1062, anoymous_9_n1216, anoymous_9_n1395);
	nor gate_anoymous_9_n198 (anoymous_9_n198, anoymous_9_n1215, anoymous_9_n1395);
	nor gate_anoymous_9_n1061 (anoymous_9_n1061, anoymous_9_n1214, anoymous_9_n1395);
	nor gate_anoymous_9_n176 (anoymous_9_n176, anoymous_9_n1213, anoymous_9_n1395);
	nor gate_anoymous_9_n1060 (anoymous_9_n1060, anoymous_9_n1212, anoymous_9_n1395);
	and gate_anoymous_9_n753 (anoymous_9_n753, anoymous_9_n1193, anoymous_9_n1209);
	xor gate_anoymous_9_n754 (anoymous_9_n754, anoymous_9_n1209, anoymous_9_n1193);
	xor gate_anoymous_9_n750 (anoymous_9_n750, anoymous_9_n1208, anoymous_9_n1192);
	and gate_anoymous_9_n749 (anoymous_9_n749, anoymous_9_n1192, anoymous_9_n1208);
	and gate_anoymous_9_n748 (anoymous_9_n748, anoymous_9_n750, anoymous_9_n1176);
	or gate_anoymous_9_n751 (anoymous_9_n751, anoymous_9_n749, anoymous_9_n748);
	xor gate_anoymous_9_n752 (anoymous_9_n752, anoymous_9_n1176, anoymous_9_n750);
	and gate_anoymous_9_n746 (anoymous_9_n746, anoymous_9_n1057, anoymous_9_n1207);
	xor gate_anoymous_9_n747 (anoymous_9_n747, anoymous_9_n1207, anoymous_9_n1057);
	xor gate_anoymous_9_n743 (anoymous_9_n743, anoymous_9_n1191, anoymous_9_n1175);
	and gate_anoymous_9_n742 (anoymous_9_n742, anoymous_9_n1175, anoymous_9_n1191);
	and gate_anoymous_9_n741 (anoymous_9_n741, anoymous_9_n747, anoymous_9_n743);
	or gate_anoymous_9_n744 (anoymous_9_n744, anoymous_9_n742, anoymous_9_n741);
	xor gate_anoymous_9_n745 (anoymous_9_n745, anoymous_9_n743, anoymous_9_n747);
	xor gate_anoymous_9_n738 (anoymous_9_n738, anoymous_9_n1206, anoymous_9_n1190);
	and gate_anoymous_9_n737 (anoymous_9_n737, anoymous_9_n1190, anoymous_9_n1206);
	and gate_anoymous_9_n736 (anoymous_9_n736, anoymous_9_n738, anoymous_9_n1174);
	or gate_anoymous_9_n739 (anoymous_9_n739, anoymous_9_n737, anoymous_9_n736);
	xor gate_anoymous_9_n740 (anoymous_9_n740, anoymous_9_n1174, anoymous_9_n738);
	xor gate_anoymous_9_n733 (anoymous_9_n733, anoymous_9_n1158, anoymous_9_n746);
	and gate_anoymous_9_n732 (anoymous_9_n732, anoymous_9_n746, anoymous_9_n1158);
	and gate_anoymous_9_n731 (anoymous_9_n731, anoymous_9_n744, anoymous_9_n733);
	or gate_anoymous_9_n734 (anoymous_9_n734, anoymous_9_n732, anoymous_9_n731);
	xor gate_anoymous_9_n735 (anoymous_9_n735, anoymous_9_n733, anoymous_9_n744);
	and gate_anoymous_9_n729 (anoymous_9_n729, anoymous_9_n1056, anoymous_9_n1205);
	xor gate_anoymous_9_n730 (anoymous_9_n730, anoymous_9_n1205, anoymous_9_n1056);
	xor gate_anoymous_9_n726 (anoymous_9_n726, anoymous_9_n1189, anoymous_9_n1173);
	and gate_anoymous_9_n725 (anoymous_9_n725, anoymous_9_n1173, anoymous_9_n1189);
	and gate_anoymous_9_n724 (anoymous_9_n724, anoymous_9_n726, anoymous_9_n1157);
	or gate_anoymous_9_n727 (anoymous_9_n727, anoymous_9_n725, anoymous_9_n724);
	xor gate_anoymous_9_n728 (anoymous_9_n728, anoymous_9_n1157, anoymous_9_n726);
	xor gate_anoymous_9_n721 (anoymous_9_n721, anoymous_9_n730, anoymous_9_n739);
	and gate_anoymous_9_n720 (anoymous_9_n720, anoymous_9_n739, anoymous_9_n730);
	and gate_anoymous_9_n719 (anoymous_9_n719, anoymous_9_n721, anoymous_9_n728);
	or gate_anoymous_9_n722 (anoymous_9_n722, anoymous_9_n720, anoymous_9_n719);
	xor gate_anoymous_9_n723 (anoymous_9_n723, anoymous_9_n728, anoymous_9_n721);
	xor gate_anoymous_9_n716 (anoymous_9_n716, anoymous_9_n1204, anoymous_9_n1188);
	and gate_anoymous_9_n715 (anoymous_9_n715, anoymous_9_n1188, anoymous_9_n1204);
	and gate_anoymous_9_n714 (anoymous_9_n714, anoymous_9_n716, anoymous_9_n1172);
	or gate_anoymous_9_n717 (anoymous_9_n717, anoymous_9_n715, anoymous_9_n714);
	xor gate_anoymous_9_n718 (anoymous_9_n718, anoymous_9_n1172, anoymous_9_n716);
	xor gate_anoymous_9_n711 (anoymous_9_n711, anoymous_9_n1156, anoymous_9_n1140);
	and gate_anoymous_9_n710 (anoymous_9_n710, anoymous_9_n1140, anoymous_9_n1156);
	and gate_anoymous_9_n709 (anoymous_9_n709, anoymous_9_n711, anoymous_9_n729);
	or gate_anoymous_9_n712 (anoymous_9_n712, anoymous_9_n710, anoymous_9_n709);
	xor gate_anoymous_9_n713 (anoymous_9_n713, anoymous_9_n729, anoymous_9_n711);
	xor gate_anoymous_9_n706 (anoymous_9_n706, anoymous_9_n727, anoymous_9_n718);
	and gate_anoymous_9_n705 (anoymous_9_n705, anoymous_9_n718, anoymous_9_n727);
	and gate_anoymous_9_n704 (anoymous_9_n704, anoymous_9_n706, anoymous_9_n713);
	or gate_anoymous_9_n707 (anoymous_9_n707, anoymous_9_n705, anoymous_9_n704);
	xor gate_anoymous_9_n708 (anoymous_9_n708, anoymous_9_n713, anoymous_9_n706);
	and gate_anoymous_9_n702 (anoymous_9_n702, anoymous_9_n1055, anoymous_9_n1203);
	xor gate_anoymous_9_n703 (anoymous_9_n703, anoymous_9_n1203, anoymous_9_n1055);
	xor gate_anoymous_9_n699 (anoymous_9_n699, anoymous_9_n1155, anoymous_9_n1187);
	and gate_anoymous_9_n698 (anoymous_9_n698, anoymous_9_n1187, anoymous_9_n1155);
	and gate_anoymous_9_n697 (anoymous_9_n697, anoymous_9_n699, anoymous_9_n1171);
	or gate_anoymous_9_n700 (anoymous_9_n700, anoymous_9_n698, anoymous_9_n697);
	xor gate_anoymous_9_n701 (anoymous_9_n701, anoymous_9_n1171, anoymous_9_n699);
	xor gate_anoymous_9_n694 (anoymous_9_n694, anoymous_9_n1139, anoymous_9_n703);
	and gate_anoymous_9_n693 (anoymous_9_n693, anoymous_9_n703, anoymous_9_n1139);
	and gate_anoymous_9_n692 (anoymous_9_n692, anoymous_9_n694, anoymous_9_n717);
	or gate_anoymous_9_n695 (anoymous_9_n695, anoymous_9_n693, anoymous_9_n692);
	xor gate_anoymous_9_n696 (anoymous_9_n696, anoymous_9_n717, anoymous_9_n694);
	xor gate_anoymous_9_n689 (anoymous_9_n689, anoymous_9_n712, anoymous_9_n701);
	and gate_anoymous_9_n688 (anoymous_9_n688, anoymous_9_n701, anoymous_9_n712);
	and gate_anoymous_9_n687 (anoymous_9_n687, anoymous_9_n696, anoymous_9_n689);
	or gate_anoymous_9_n690 (anoymous_9_n690, anoymous_9_n688, anoymous_9_n687);
	xor gate_anoymous_9_n691 (anoymous_9_n691, anoymous_9_n689, anoymous_9_n696);
	xor gate_anoymous_9_n684 (anoymous_9_n684, anoymous_9_n1202, anoymous_9_n1186);
	and gate_anoymous_9_n683 (anoymous_9_n683, anoymous_9_n1186, anoymous_9_n1202);
	and gate_anoymous_9_n682 (anoymous_9_n682, anoymous_9_n684, anoymous_9_n1170);
	or gate_anoymous_9_n685 (anoymous_9_n685, anoymous_9_n683, anoymous_9_n682);
	xor gate_anoymous_9_n686 (anoymous_9_n686, anoymous_9_n1170, anoymous_9_n684);
	xor gate_anoymous_9_n679 (anoymous_9_n679, anoymous_9_n1154, anoymous_9_n1138);
	and gate_anoymous_9_n678 (anoymous_9_n678, anoymous_9_n1138, anoymous_9_n1154);
	and gate_anoymous_9_n677 (anoymous_9_n677, anoymous_9_n679, anoymous_9_n1122);
	or gate_anoymous_9_n680 (anoymous_9_n680, anoymous_9_n678, anoymous_9_n677);
	xor gate_anoymous_9_n681 (anoymous_9_n681, anoymous_9_n1122, anoymous_9_n679);
	xor gate_anoymous_9_n674 (anoymous_9_n674, anoymous_9_n702, anoymous_9_n700);
	and gate_anoymous_9_n673 (anoymous_9_n673, anoymous_9_n700, anoymous_9_n702);
	and gate_anoymous_9_n672 (anoymous_9_n672, anoymous_9_n674, anoymous_9_n686);
	or gate_anoymous_9_n675 (anoymous_9_n675, anoymous_9_n673, anoymous_9_n672);
	xor gate_anoymous_9_n676 (anoymous_9_n676, anoymous_9_n686, anoymous_9_n674);
	xor gate_anoymous_9_n669 (anoymous_9_n669, anoymous_9_n681, anoymous_9_n695);
	and gate_anoymous_9_n668 (anoymous_9_n668, anoymous_9_n695, anoymous_9_n681);
	and gate_anoymous_9_n667 (anoymous_9_n667, anoymous_9_n676, anoymous_9_n669);
	or gate_anoymous_9_n670 (anoymous_9_n670, anoymous_9_n668, anoymous_9_n667);
	xor gate_anoymous_9_n671 (anoymous_9_n671, anoymous_9_n669, anoymous_9_n676);
	and gate_anoymous_9_n665 (anoymous_9_n665, anoymous_9_n1054, anoymous_9_n1201);
	xor gate_anoymous_9_n666 (anoymous_9_n666, anoymous_9_n1201, anoymous_9_n1054);
	xor gate_anoymous_9_n662 (anoymous_9_n662, anoymous_9_n1153, anoymous_9_n1137);
	and gate_anoymous_9_n661 (anoymous_9_n661, anoymous_9_n1137, anoymous_9_n1153);
	and gate_anoymous_9_n660 (anoymous_9_n660, anoymous_9_n662, anoymous_9_n1121);
	or gate_anoymous_9_n663 (anoymous_9_n663, anoymous_9_n661, anoymous_9_n660);
	xor gate_anoymous_9_n664 (anoymous_9_n664, anoymous_9_n1121, anoymous_9_n662);
	xor gate_anoymous_9_n657 (anoymous_9_n657, anoymous_9_n1185, anoymous_9_n1169);
	and gate_anoymous_9_n656 (anoymous_9_n656, anoymous_9_n1169, anoymous_9_n1185);
	and gate_anoymous_9_n655 (anoymous_9_n655, anoymous_9_n666, anoymous_9_n657);
	or gate_anoymous_9_n658 (anoymous_9_n658, anoymous_9_n656, anoymous_9_n655);
	xor gate_anoymous_9_n659 (anoymous_9_n659, anoymous_9_n657, anoymous_9_n666);
	xor gate_anoymous_9_n652 (anoymous_9_n652, anoymous_9_n685, anoymous_9_n680);
	and gate_anoymous_9_n651 (anoymous_9_n651, anoymous_9_n680, anoymous_9_n685);
	and gate_anoymous_9_n650 (anoymous_9_n650, anoymous_9_n652, anoymous_9_n664);
	or gate_anoymous_9_n653 (anoymous_9_n653, anoymous_9_n651, anoymous_9_n650);
	xor gate_anoymous_9_n654 (anoymous_9_n654, anoymous_9_n664, anoymous_9_n652);
	xor gate_anoymous_9_n647 (anoymous_9_n647, anoymous_9_n659, anoymous_9_n675);
	and gate_anoymous_9_n646 (anoymous_9_n646, anoymous_9_n675, anoymous_9_n659);
	and gate_anoymous_9_n645 (anoymous_9_n645, anoymous_9_n647, anoymous_9_n654);
	or gate_anoymous_9_n648 (anoymous_9_n648, anoymous_9_n646, anoymous_9_n645);
	xor gate_anoymous_9_n649 (anoymous_9_n649, anoymous_9_n654, anoymous_9_n647);
	xor gate_anoymous_9_n642 (anoymous_9_n642, anoymous_9_n1200, anoymous_9_n1184);
	and gate_anoymous_9_n641 (anoymous_9_n641, anoymous_9_n1184, anoymous_9_n1200);
	and gate_anoymous_9_n640 (anoymous_9_n640, anoymous_9_n642, anoymous_9_n1168);
	or gate_anoymous_9_n643 (anoymous_9_n643, anoymous_9_n641, anoymous_9_n640);
	xor gate_anoymous_9_n644 (anoymous_9_n644, anoymous_9_n1168, anoymous_9_n642);
	xor gate_anoymous_9_n637 (anoymous_9_n637, anoymous_9_n1152, anoymous_9_n1136);
	and gate_anoymous_9_n636 (anoymous_9_n636, anoymous_9_n1136, anoymous_9_n1152);
	and gate_anoymous_9_n635 (anoymous_9_n635, anoymous_9_n637, anoymous_9_n1120);
	or gate_anoymous_9_n638 (anoymous_9_n638, anoymous_9_n636, anoymous_9_n635);
	xor gate_anoymous_9_n639 (anoymous_9_n639, anoymous_9_n1120, anoymous_9_n637);
	xor gate_anoymous_9_n632 (anoymous_9_n632, anoymous_9_n1104, anoymous_9_n665);
	and gate_anoymous_9_n631 (anoymous_9_n631, anoymous_9_n665, anoymous_9_n1104);
	and gate_anoymous_9_n630 (anoymous_9_n630, anoymous_9_n663, anoymous_9_n632);
	or gate_anoymous_9_n633 (anoymous_9_n633, anoymous_9_n631, anoymous_9_n630);
	xor gate_anoymous_9_n634 (anoymous_9_n634, anoymous_9_n632, anoymous_9_n663);
	xor gate_anoymous_9_n627 (anoymous_9_n627, anoymous_9_n658, anoymous_9_n644);
	and gate_anoymous_9_n626 (anoymous_9_n626, anoymous_9_n644, anoymous_9_n658);
	and gate_anoymous_9_n625 (anoymous_9_n625, anoymous_9_n627, anoymous_9_n639);
	or gate_anoymous_9_n628 (anoymous_9_n628, anoymous_9_n626, anoymous_9_n625);
	xor gate_anoymous_9_n629 (anoymous_9_n629, anoymous_9_n639, anoymous_9_n627);
	xor gate_anoymous_9_n622 (anoymous_9_n622, anoymous_9_n634, anoymous_9_n653);
	and gate_anoymous_9_n621 (anoymous_9_n621, anoymous_9_n653, anoymous_9_n634);
	and gate_anoymous_9_n620 (anoymous_9_n620, anoymous_9_n622, anoymous_9_n629);
	or gate_anoymous_9_n623 (anoymous_9_n623, anoymous_9_n621, anoymous_9_n620);
	xor gate_anoymous_9_n624 (anoymous_9_n624, anoymous_9_n629, anoymous_9_n622);
	and gate_anoymous_9_n618 (anoymous_9_n618, anoymous_9_n1053, anoymous_9_n1199);
	xor gate_anoymous_9_n619 (anoymous_9_n619, anoymous_9_n1199, anoymous_9_n1053);
	xor gate_anoymous_9_n615 (anoymous_9_n615, anoymous_9_n1135, anoymous_9_n1151);
	and gate_anoymous_9_n614 (anoymous_9_n614, anoymous_9_n1151, anoymous_9_n1135);
	and gate_anoymous_9_n613 (anoymous_9_n613, anoymous_9_n615, anoymous_9_n1119);
	or gate_anoymous_9_n616 (anoymous_9_n616, anoymous_9_n614, anoymous_9_n613);
	xor gate_anoymous_9_n617 (anoymous_9_n617, anoymous_9_n1119, anoymous_9_n615);
	xor gate_anoymous_9_n610 (anoymous_9_n610, anoymous_9_n1183, anoymous_9_n1167);
	and gate_anoymous_9_n609 (anoymous_9_n609, anoymous_9_n1167, anoymous_9_n1183);
	and gate_anoymous_9_n608 (anoymous_9_n608, anoymous_9_n610, anoymous_9_n1103);
	or gate_anoymous_9_n611 (anoymous_9_n611, anoymous_9_n609, anoymous_9_n608);
	xor gate_anoymous_9_n612 (anoymous_9_n612, anoymous_9_n1103, anoymous_9_n610);
	xor gate_anoymous_9_n605 (anoymous_9_n605, anoymous_9_n619, anoymous_9_n643);
	and gate_anoymous_9_n604 (anoymous_9_n604, anoymous_9_n643, anoymous_9_n619);
	and gate_anoymous_9_n603 (anoymous_9_n603, anoymous_9_n605, anoymous_9_n638);
	or gate_anoymous_9_n606 (anoymous_9_n606, anoymous_9_n604, anoymous_9_n603);
	xor gate_anoymous_9_n607 (anoymous_9_n607, anoymous_9_n638, anoymous_9_n605);
	xor gate_anoymous_9_n600 (anoymous_9_n600, anoymous_9_n612, anoymous_9_n617);
	and gate_anoymous_9_n599 (anoymous_9_n599, anoymous_9_n617, anoymous_9_n612);
	and gate_anoymous_9_n598 (anoymous_9_n598, anoymous_9_n600, anoymous_9_n633);
	or gate_anoymous_9_n601 (anoymous_9_n601, anoymous_9_n599, anoymous_9_n598);
	xor gate_anoymous_9_n602 (anoymous_9_n602, anoymous_9_n633, anoymous_9_n600);
	xor gate_anoymous_9_n595 (anoymous_9_n595, anoymous_9_n607, anoymous_9_n628);
	and gate_anoymous_9_n594 (anoymous_9_n594, anoymous_9_n628, anoymous_9_n607);
	and gate_anoymous_9_n593 (anoymous_9_n593, anoymous_9_n595, anoymous_9_n602);
	or gate_anoymous_9_n596 (anoymous_9_n596, anoymous_9_n594, anoymous_9_n593);
	xor gate_anoymous_9_n597 (anoymous_9_n597, anoymous_9_n602, anoymous_9_n595);
	xor gate_anoymous_9_n590 (anoymous_9_n590, anoymous_9_n1198, anoymous_9_n1182);
	and gate_anoymous_9_n589 (anoymous_9_n589, anoymous_9_n1182, anoymous_9_n1198);
	and gate_anoymous_9_n588 (anoymous_9_n588, anoymous_9_n590, anoymous_9_n1166);
	or gate_anoymous_9_n591 (anoymous_9_n591, anoymous_9_n589, anoymous_9_n588);
	xor gate_anoymous_9_n592 (anoymous_9_n592, anoymous_9_n1166, anoymous_9_n590);
	xor gate_anoymous_9_n585 (anoymous_9_n585, anoymous_9_n1150, anoymous_9_n1134);
	and gate_anoymous_9_n584 (anoymous_9_n584, anoymous_9_n1134, anoymous_9_n1150);
	and gate_anoymous_9_n583 (anoymous_9_n583, anoymous_9_n585, anoymous_9_n1118);
	or gate_anoymous_9_n586 (anoymous_9_n586, anoymous_9_n584, anoymous_9_n583);
	xor gate_anoymous_9_n587 (anoymous_9_n587, anoymous_9_n1118, anoymous_9_n585);
	xor gate_anoymous_9_n580 (anoymous_9_n580, anoymous_9_n1102, anoymous_9_n1086);
	and gate_anoymous_9_n579 (anoymous_9_n579, anoymous_9_n1086, anoymous_9_n1102);
	and gate_anoymous_9_n578 (anoymous_9_n578, anoymous_9_n580, anoymous_9_n618);
	or gate_anoymous_9_n581 (anoymous_9_n581, anoymous_9_n579, anoymous_9_n578);
	xor gate_anoymous_9_n582 (anoymous_9_n582, anoymous_9_n618, anoymous_9_n580);
	xor gate_anoymous_9_n575 (anoymous_9_n575, anoymous_9_n616, anoymous_9_n611);
	and gate_anoymous_9_n574 (anoymous_9_n574, anoymous_9_n611, anoymous_9_n616);
	and gate_anoymous_9_n573 (anoymous_9_n573, anoymous_9_n575, anoymous_9_n592);
	or gate_anoymous_9_n576 (anoymous_9_n576, anoymous_9_n574, anoymous_9_n573);
	xor gate_anoymous_9_n577 (anoymous_9_n577, anoymous_9_n592, anoymous_9_n575);
	xor gate_anoymous_9_n570 (anoymous_9_n570, anoymous_9_n587, anoymous_9_n582);
	and gate_anoymous_9_n569 (anoymous_9_n569, anoymous_9_n582, anoymous_9_n587);
	and gate_anoymous_9_n568 (anoymous_9_n568, anoymous_9_n606, anoymous_9_n570);
	or gate_anoymous_9_n571 (anoymous_9_n571, anoymous_9_n569, anoymous_9_n568);
	xor gate_anoymous_9_n572 (anoymous_9_n572, anoymous_9_n570, anoymous_9_n606);
	xor gate_anoymous_9_n565 (anoymous_9_n565, anoymous_9_n577, anoymous_9_n601);
	and gate_anoymous_9_n564 (anoymous_9_n564, anoymous_9_n601, anoymous_9_n577);
	and gate_anoymous_9_n563 (anoymous_9_n563, anoymous_9_n565, anoymous_9_n572);
	or gate_anoymous_9_n566 (anoymous_9_n566, anoymous_9_n564, anoymous_9_n563);
	xor gate_anoymous_9_n567 (anoymous_9_n567, anoymous_9_n572, anoymous_9_n565);
	and gate_anoymous_9_n561 (anoymous_9_n561, anoymous_9_n1052, anoymous_9_n1197);
	xor gate_anoymous_9_n562 (anoymous_9_n562, anoymous_9_n1197, anoymous_9_n1052);
	xor gate_anoymous_9_n558 (anoymous_9_n558, anoymous_9_n1133, anoymous_9_n1117);
	and gate_anoymous_9_n557 (anoymous_9_n557, anoymous_9_n1117, anoymous_9_n1133);
	and gate_anoymous_9_n556 (anoymous_9_n556, anoymous_9_n558, anoymous_9_n1101);
	or gate_anoymous_9_n559 (anoymous_9_n559, anoymous_9_n557, anoymous_9_n556);
	xor gate_anoymous_9_n560 (anoymous_9_n560, anoymous_9_n1101, anoymous_9_n558);
	xor gate_anoymous_9_n553 (anoymous_9_n553, anoymous_9_n1085, anoymous_9_n1149);
	and gate_anoymous_9_n552 (anoymous_9_n552, anoymous_9_n1149, anoymous_9_n1085);
	and gate_anoymous_9_n551 (anoymous_9_n551, anoymous_9_n553, anoymous_9_n1181);
	or gate_anoymous_9_n554 (anoymous_9_n554, anoymous_9_n552, anoymous_9_n551);
	xor gate_anoymous_9_n555 (anoymous_9_n555, anoymous_9_n1181, anoymous_9_n553);
	xor gate_anoymous_9_n548 (anoymous_9_n548, anoymous_9_n1165, anoymous_9_n562);
	and gate_anoymous_9_n547 (anoymous_9_n547, anoymous_9_n562, anoymous_9_n1165);
	and gate_anoymous_9_n546 (anoymous_9_n546, anoymous_9_n548, anoymous_9_n591);
	or gate_anoymous_9_n549 (anoymous_9_n549, anoymous_9_n547, anoymous_9_n546);
	xor gate_anoymous_9_n550 (anoymous_9_n550, anoymous_9_n591, anoymous_9_n548);
	xor gate_anoymous_9_n543 (anoymous_9_n543, anoymous_9_n586, anoymous_9_n581);
	and gate_anoymous_9_n542 (anoymous_9_n542, anoymous_9_n581, anoymous_9_n586);
	and gate_anoymous_9_n541 (anoymous_9_n541, anoymous_9_n543, anoymous_9_n555);
	or gate_anoymous_9_n544 (anoymous_9_n544, anoymous_9_n542, anoymous_9_n541);
	xor gate_anoymous_9_n545 (anoymous_9_n545, anoymous_9_n555, anoymous_9_n543);
	xor gate_anoymous_9_n538 (anoymous_9_n538, anoymous_9_n560, anoymous_9_n550);
	and gate_anoymous_9_n537 (anoymous_9_n537, anoymous_9_n550, anoymous_9_n560);
	and gate_anoymous_9_n536 (anoymous_9_n536, anoymous_9_n538, anoymous_9_n576);
	or gate_anoymous_9_n539 (anoymous_9_n539, anoymous_9_n537, anoymous_9_n536);
	xor gate_anoymous_9_n540 (anoymous_9_n540, anoymous_9_n576, anoymous_9_n538);
	xor gate_anoymous_9_n533 (anoymous_9_n533, anoymous_9_n545, anoymous_9_n571);
	and gate_anoymous_9_n532 (anoymous_9_n532, anoymous_9_n571, anoymous_9_n545);
	and gate_anoymous_9_n531 (anoymous_9_n531, anoymous_9_n540, anoymous_9_n533);
	or gate_anoymous_9_n534 (anoymous_9_n534, anoymous_9_n532, anoymous_9_n531);
	xor gate_anoymous_9_n535 (anoymous_9_n535, anoymous_9_n533, anoymous_9_n540);
	xor gate_anoymous_9_n528 (anoymous_9_n528, anoymous_9_n1068, anoymous_9_n1196);
	and gate_anoymous_9_n527 (anoymous_9_n527, anoymous_9_n1196, anoymous_9_n1068);
	and gate_anoymous_9_n526 (anoymous_9_n526, anoymous_9_n528, anoymous_9_n1180);
	or gate_anoymous_9_n529 (anoymous_9_n529, anoymous_9_n527, anoymous_9_n526);
	xor gate_anoymous_9_n530 (anoymous_9_n530, anoymous_9_n1180, anoymous_9_n528);
	xor gate_anoymous_9_n523 (anoymous_9_n523, anoymous_9_n1164, anoymous_9_n1148);
	and gate_anoymous_9_n522 (anoymous_9_n522, anoymous_9_n1148, anoymous_9_n1164);
	and gate_anoymous_9_n521 (anoymous_9_n521, anoymous_9_n523, anoymous_9_n1132);
	or gate_anoymous_9_n524 (anoymous_9_n524, anoymous_9_n522, anoymous_9_n521);
	xor gate_anoymous_9_n525 (anoymous_9_n525, anoymous_9_n1132, anoymous_9_n523);
	xor gate_anoymous_9_n518 (anoymous_9_n518, anoymous_9_n1116, anoymous_9_n1100);
	and gate_anoymous_9_n517 (anoymous_9_n517, anoymous_9_n1100, anoymous_9_n1116);
	and gate_anoymous_9_n516 (anoymous_9_n516, anoymous_9_n518, anoymous_9_n1084);
	or gate_anoymous_9_n519 (anoymous_9_n519, anoymous_9_n517, anoymous_9_n516);
	xor gate_anoymous_9_n520 (anoymous_9_n520, anoymous_9_n1084, anoymous_9_n518);
	xor gate_anoymous_9_n513 (anoymous_9_n513, anoymous_9_n561, anoymous_9_n559);
	and gate_anoymous_9_n512 (anoymous_9_n512, anoymous_9_n559, anoymous_9_n561);
	and gate_anoymous_9_n511 (anoymous_9_n511, anoymous_9_n513, anoymous_9_n554);
	or gate_anoymous_9_n514 (anoymous_9_n514, anoymous_9_n512, anoymous_9_n511);
	xor gate_anoymous_9_n515 (anoymous_9_n515, anoymous_9_n554, anoymous_9_n513);
	xor gate_anoymous_9_n508 (anoymous_9_n508, anoymous_9_n530, anoymous_9_n520);
	and gate_anoymous_9_n507 (anoymous_9_n507, anoymous_9_n520, anoymous_9_n530);
	and gate_anoymous_9_n506 (anoymous_9_n506, anoymous_9_n508, anoymous_9_n525);
	or gate_anoymous_9_n509 (anoymous_9_n509, anoymous_9_n507, anoymous_9_n506);
	xor gate_anoymous_9_n510 (anoymous_9_n510, anoymous_9_n525, anoymous_9_n508);
	xor gate_anoymous_9_n503 (anoymous_9_n503, anoymous_9_n549, anoymous_9_n544);
	and gate_anoymous_9_n502 (anoymous_9_n502, anoymous_9_n544, anoymous_9_n549);
	and gate_anoymous_9_n501 (anoymous_9_n501, anoymous_9_n503, anoymous_9_n515);
	or gate_anoymous_9_n504 (anoymous_9_n504, anoymous_9_n502, anoymous_9_n501);
	xor gate_anoymous_9_n505 (anoymous_9_n505, anoymous_9_n515, anoymous_9_n503);
	xor gate_anoymous_9_n498 (anoymous_9_n498, anoymous_9_n510, anoymous_9_n539);
	and gate_anoymous_9_n497 (anoymous_9_n497, anoymous_9_n539, anoymous_9_n510);
	and gate_anoymous_9_n496 (anoymous_9_n496, anoymous_9_n498, anoymous_9_n505);
	or gate_anoymous_9_n499 (anoymous_9_n499, anoymous_9_n497, anoymous_9_n496);
	xor gate_anoymous_9_n500 (anoymous_9_n500, anoymous_9_n505, anoymous_9_n498);
	not gate_anoymous_9_n495 (anoymous_9_n495, anoymous_9_n458);
	xor gate_anoymous_9_n492 (anoymous_9_n492, anoymous_9_n495, anoymous_9_n1099);
	and gate_anoymous_9_n491 (anoymous_9_n491, anoymous_9_n1099, anoymous_9_n495);
	and gate_anoymous_9_n490 (anoymous_9_n490, anoymous_9_n492, anoymous_9_n1147);
	or gate_anoymous_9_n493 (anoymous_9_n493, anoymous_9_n491, anoymous_9_n490);
	xor gate_anoymous_9_n494 (anoymous_9_n494, anoymous_9_n1147, anoymous_9_n492);
	xor gate_anoymous_9_n487 (anoymous_9_n487, anoymous_9_n1131, anoymous_9_n1163);
	and gate_anoymous_9_n486 (anoymous_9_n486, anoymous_9_n1163, anoymous_9_n1131);
	and gate_anoymous_9_n485 (anoymous_9_n485, anoymous_9_n487, anoymous_9_n1115);
	or gate_anoymous_9_n488 (anoymous_9_n488, anoymous_9_n486, anoymous_9_n485);
	xor gate_anoymous_9_n489 (anoymous_9_n489, anoymous_9_n1115, anoymous_9_n487);
	xor gate_anoymous_9_n482 (anoymous_9_n482, anoymous_9_n1179, anoymous_9_n1083);
	and gate_anoymous_9_n481 (anoymous_9_n481, anoymous_9_n1083, anoymous_9_n1179);
	and gate_anoymous_9_n480 (anoymous_9_n480, anoymous_9_n482, anoymous_9_n1195);
	or gate_anoymous_9_n483 (anoymous_9_n483, anoymous_9_n481, anoymous_9_n480);
	xor gate_anoymous_9_n484 (anoymous_9_n484, anoymous_9_n1195, anoymous_9_n482);
	xor gate_anoymous_9_n477 (anoymous_9_n477, anoymous_9_n529, anoymous_9_n524);
	and gate_anoymous_9_n476 (anoymous_9_n476, anoymous_9_n524, anoymous_9_n529);
	and gate_anoymous_9_n475 (anoymous_9_n475, anoymous_9_n477, anoymous_9_n519);
	or gate_anoymous_9_n478 (anoymous_9_n478, anoymous_9_n476, anoymous_9_n475);
	xor gate_anoymous_9_n479 (anoymous_9_n479, anoymous_9_n519, anoymous_9_n477);
	xor gate_anoymous_9_n472 (anoymous_9_n472, anoymous_9_n494, anoymous_9_n484);
	and gate_anoymous_9_n471 (anoymous_9_n471, anoymous_9_n484, anoymous_9_n494);
	and gate_anoymous_9_n470 (anoymous_9_n470, anoymous_9_n472, anoymous_9_n489);
	or gate_anoymous_9_n473 (anoymous_9_n473, anoymous_9_n471, anoymous_9_n470);
	xor gate_anoymous_9_n474 (anoymous_9_n474, anoymous_9_n489, anoymous_9_n472);
	xor gate_anoymous_9_n467 (anoymous_9_n467, anoymous_9_n514, anoymous_9_n479);
	and gate_anoymous_9_n466 (anoymous_9_n466, anoymous_9_n479, anoymous_9_n514);
	and gate_anoymous_9_n465 (anoymous_9_n465, anoymous_9_n467, anoymous_9_n509);
	or gate_anoymous_9_n468 (anoymous_9_n468, anoymous_9_n466, anoymous_9_n465);
	xor gate_anoymous_9_n469 (anoymous_9_n469, anoymous_9_n509, anoymous_9_n467);
	xor gate_anoymous_9_n462 (anoymous_9_n462, anoymous_9_n474, anoymous_9_n504);
	and gate_anoymous_9_n461 (anoymous_9_n461, anoymous_9_n504, anoymous_9_n474);
	and gate_anoymous_9_n460 (anoymous_9_n460, anoymous_9_n462, anoymous_9_n469);
	or gate_anoymous_9_n463 (anoymous_9_n463, anoymous_9_n461, anoymous_9_n460);
	xor gate_anoymous_9_n464 (anoymous_9_n464, anoymous_9_n469, anoymous_9_n462);
	not gate_anoymous_9_n459 (anoymous_9_n459, anoymous_9_n458);
	xor gate_anoymous_9_n455 (anoymous_9_n455, anoymous_9_n1067, anoymous_9_n459);
	and gate_anoymous_9_n454 (anoymous_9_n454, anoymous_9_n459, anoymous_9_n1067);
	and gate_anoymous_9_n453 (anoymous_9_n453, anoymous_9_n455, anoymous_9_n1178);
	or gate_anoymous_9_n456 (anoymous_9_n456, anoymous_9_n454, anoymous_9_n453);
	xor gate_anoymous_9_n457 (anoymous_9_n457, anoymous_9_n1178, anoymous_9_n455);
	xor gate_anoymous_9_n450 (anoymous_9_n450, anoymous_9_n1114, anoymous_9_n1098);
	and gate_anoymous_9_n449 (anoymous_9_n449, anoymous_9_n1098, anoymous_9_n1114);
	and gate_anoymous_9_n448 (anoymous_9_n448, anoymous_9_n450, anoymous_9_n1130);
	or gate_anoymous_9_n451 (anoymous_9_n451, anoymous_9_n449, anoymous_9_n448);
	xor gate_anoymous_9_n452 (anoymous_9_n452, anoymous_9_n1130, anoymous_9_n450);
	xor gate_anoymous_9_n445 (anoymous_9_n445, anoymous_9_n1162, anoymous_9_n1146);
	and gate_anoymous_9_n444 (anoymous_9_n444, anoymous_9_n1146, anoymous_9_n1162);
	and gate_anoymous_9_n443 (anoymous_9_n443, anoymous_9_n445, anoymous_9_n1082);
	or gate_anoymous_9_n446 (anoymous_9_n446, anoymous_9_n444, anoymous_9_n443);
	xor gate_anoymous_9_n447 (anoymous_9_n447, anoymous_9_n1082, anoymous_9_n445);
	xor gate_anoymous_9_n440 (anoymous_9_n440, anoymous_9_n457, anoymous_9_n493);
	and gate_anoymous_9_n439 (anoymous_9_n439, anoymous_9_n493, anoymous_9_n457);
	and gate_anoymous_9_n438 (anoymous_9_n438, anoymous_9_n440, anoymous_9_n488);
	or gate_anoymous_9_n441 (anoymous_9_n441, anoymous_9_n439, anoymous_9_n438);
	xor gate_anoymous_9_n442 (anoymous_9_n442, anoymous_9_n488, anoymous_9_n440);
	xor gate_anoymous_9_n435 (anoymous_9_n435, anoymous_9_n483, anoymous_9_n447);
	and gate_anoymous_9_n434 (anoymous_9_n434, anoymous_9_n447, anoymous_9_n483);
	and gate_anoymous_9_n433 (anoymous_9_n433, anoymous_9_n435, anoymous_9_n452);
	or gate_anoymous_9_n436 (anoymous_9_n436, anoymous_9_n434, anoymous_9_n433);
	xor gate_anoymous_9_n437 (anoymous_9_n437, anoymous_9_n452, anoymous_9_n435);
	xor gate_anoymous_9_n430 (anoymous_9_n430, anoymous_9_n478, anoymous_9_n442);
	and gate_anoymous_9_n429 (anoymous_9_n429, anoymous_9_n442, anoymous_9_n478);
	and gate_anoymous_9_n428 (anoymous_9_n428, anoymous_9_n430, anoymous_9_n473);
	or gate_anoymous_9_n431 (anoymous_9_n431, anoymous_9_n429, anoymous_9_n428);
	xor gate_anoymous_9_n432 (anoymous_9_n432, anoymous_9_n473, anoymous_9_n430);
	xor gate_anoymous_9_n425 (anoymous_9_n425, anoymous_9_n437, anoymous_9_n468);
	and gate_anoymous_9_n424 (anoymous_9_n424, anoymous_9_n468, anoymous_9_n437);
	and gate_anoymous_9_n423 (anoymous_9_n423, anoymous_9_n425, anoymous_9_n432);
	or gate_anoymous_9_n426 (anoymous_9_n426, anoymous_9_n424, anoymous_9_n423);
	xor gate_anoymous_9_n427 (anoymous_9_n427, anoymous_9_n432, anoymous_9_n425);
	xor gate_anoymous_9_n420 (anoymous_9_n420, anoymous_9_n458, anoymous_9_n1066);
	and gate_anoymous_9_n419 (anoymous_9_n419, anoymous_9_n1066, anoymous_9_n458);
	and gate_anoymous_9_n418 (anoymous_9_n418, anoymous_9_n420, anoymous_9_n1129);
	or gate_anoymous_9_n421 (anoymous_9_n421, anoymous_9_n419, anoymous_9_n418);
	xor gate_anoymous_9_n422 (anoymous_9_n422, anoymous_9_n1129, anoymous_9_n420);
	xor gate_anoymous_9_n415 (anoymous_9_n415, anoymous_9_n1113, anoymous_9_n1097);
	and gate_anoymous_9_n414 (anoymous_9_n414, anoymous_9_n1097, anoymous_9_n1113);
	and gate_anoymous_9_n413 (anoymous_9_n413, anoymous_9_n415, anoymous_9_n1145);
	or gate_anoymous_9_n416 (anoymous_9_n416, anoymous_9_n414, anoymous_9_n413);
	xor gate_anoymous_9_n417 (anoymous_9_n417, anoymous_9_n1145, anoymous_9_n415);
	xor gate_anoymous_9_n410 (anoymous_9_n410, anoymous_9_n1161, anoymous_9_n1081);
	and gate_anoymous_9_n409 (anoymous_9_n409, anoymous_9_n1081, anoymous_9_n1161);
	and gate_anoymous_9_n408 (anoymous_9_n408, anoymous_9_n410, anoymous_9_n1177);
	or gate_anoymous_9_n411 (anoymous_9_n411, anoymous_9_n409, anoymous_9_n408);
	xor gate_anoymous_9_n412 (anoymous_9_n412, anoymous_9_n1177, anoymous_9_n410);
	xor gate_anoymous_9_n405 (anoymous_9_n405, anoymous_9_n456, anoymous_9_n422);
	and gate_anoymous_9_n404 (anoymous_9_n404, anoymous_9_n422, anoymous_9_n456);
	and gate_anoymous_9_n403 (anoymous_9_n403, anoymous_9_n405, anoymous_9_n451);
	or gate_anoymous_9_n406 (anoymous_9_n406, anoymous_9_n404, anoymous_9_n403);
	xor gate_anoymous_9_n407 (anoymous_9_n407, anoymous_9_n451, anoymous_9_n405);
	xor gate_anoymous_9_n400 (anoymous_9_n400, anoymous_9_n446, anoymous_9_n412);
	and gate_anoymous_9_n399 (anoymous_9_n399, anoymous_9_n412, anoymous_9_n446);
	and gate_anoymous_9_n398 (anoymous_9_n398, anoymous_9_n400, anoymous_9_n417);
	or gate_anoymous_9_n401 (anoymous_9_n401, anoymous_9_n399, anoymous_9_n398);
	xor gate_anoymous_9_n402 (anoymous_9_n402, anoymous_9_n417, anoymous_9_n400);
	xor gate_anoymous_9_n395 (anoymous_9_n395, anoymous_9_n407, anoymous_9_n441);
	and gate_anoymous_9_n394 (anoymous_9_n394, anoymous_9_n441, anoymous_9_n407);
	and gate_anoymous_9_n393 (anoymous_9_n393, anoymous_9_n395, anoymous_9_n436);
	or gate_anoymous_9_n396 (anoymous_9_n396, anoymous_9_n394, anoymous_9_n393);
	xor gate_anoymous_9_n397 (anoymous_9_n397, anoymous_9_n436, anoymous_9_n395);
	xor gate_anoymous_9_n390 (anoymous_9_n390, anoymous_9_n402, anoymous_9_n431);
	and gate_anoymous_9_n389 (anoymous_9_n389, anoymous_9_n431, anoymous_9_n402);
	and gate_anoymous_9_n388 (anoymous_9_n388, anoymous_9_n390, anoymous_9_n397);
	or gate_anoymous_9_n391 (anoymous_9_n391, anoymous_9_n389, anoymous_9_n388);
	xor gate_anoymous_9_n392 (anoymous_9_n392, anoymous_9_n397, anoymous_9_n390);
	not gate_anoymous_9_n387 (anoymous_9_n387, anoymous_9_n386);
	xor gate_anoymous_9_n383 (anoymous_9_n383, anoymous_9_n387, anoymous_9_n1160);
	and gate_anoymous_9_n382 (anoymous_9_n382, anoymous_9_n1160, anoymous_9_n387);
	and gate_anoymous_9_n381 (anoymous_9_n381, anoymous_9_n383, anoymous_9_n1144);
	or gate_anoymous_9_n384 (anoymous_9_n384, anoymous_9_n382, anoymous_9_n381);
	xor gate_anoymous_9_n385 (anoymous_9_n385, anoymous_9_n1144, anoymous_9_n383);
	xor gate_anoymous_9_n378 (anoymous_9_n378, anoymous_9_n1128, anoymous_9_n1112);
	and gate_anoymous_9_n377 (anoymous_9_n377, anoymous_9_n1112, anoymous_9_n1128);
	and gate_anoymous_9_n376 (anoymous_9_n376, anoymous_9_n378, anoymous_9_n1080);
	or gate_anoymous_9_n379 (anoymous_9_n379, anoymous_9_n377, anoymous_9_n376);
	xor gate_anoymous_9_n380 (anoymous_9_n380, anoymous_9_n1080, anoymous_9_n378);
	xor gate_anoymous_9_n373 (anoymous_9_n373, anoymous_9_n1096, anoymous_9_n421);
	and gate_anoymous_9_n372 (anoymous_9_n372, anoymous_9_n421, anoymous_9_n1096);
	and gate_anoymous_9_n371 (anoymous_9_n371, anoymous_9_n416, anoymous_9_n373);
	or gate_anoymous_9_n374 (anoymous_9_n374, anoymous_9_n372, anoymous_9_n371);
	xor gate_anoymous_9_n375 (anoymous_9_n375, anoymous_9_n373, anoymous_9_n416);
	xor gate_anoymous_9_n368 (anoymous_9_n368, anoymous_9_n411, anoymous_9_n385);
	and gate_anoymous_9_n367 (anoymous_9_n367, anoymous_9_n385, anoymous_9_n411);
	and gate_anoymous_9_n366 (anoymous_9_n366, anoymous_9_n368, anoymous_9_n380);
	or gate_anoymous_9_n369 (anoymous_9_n369, anoymous_9_n367, anoymous_9_n366);
	xor gate_anoymous_9_n370 (anoymous_9_n370, anoymous_9_n380, anoymous_9_n368);
	xor gate_anoymous_9_n363 (anoymous_9_n363, anoymous_9_n375, anoymous_9_n406);
	and gate_anoymous_9_n362 (anoymous_9_n362, anoymous_9_n406, anoymous_9_n375);
	and gate_anoymous_9_n361 (anoymous_9_n361, anoymous_9_n363, anoymous_9_n401);
	or gate_anoymous_9_n364 (anoymous_9_n364, anoymous_9_n362, anoymous_9_n361);
	xor gate_anoymous_9_n365 (anoymous_9_n365, anoymous_9_n401, anoymous_9_n363);
	xor gate_anoymous_9_n358 (anoymous_9_n358, anoymous_9_n370, anoymous_9_n365);
	and gate_anoymous_9_n357 (anoymous_9_n357, anoymous_9_n365, anoymous_9_n370);
	and gate_anoymous_9_n356 (anoymous_9_n356, anoymous_9_n358, anoymous_9_n396);
	or gate_anoymous_9_n359 (anoymous_9_n359, anoymous_9_n357, anoymous_9_n356);
	xor gate_anoymous_9_n360 (anoymous_9_n360, anoymous_9_n396, anoymous_9_n358);
	xor gate_anoymous_9_n353 (anoymous_9_n353, anoymous_9_n386, anoymous_9_n1065);
	and gate_anoymous_9_n352 (anoymous_9_n352, anoymous_9_n1065, anoymous_9_n386);
	and gate_anoymous_9_n351 (anoymous_9_n351, anoymous_9_n353, anoymous_9_n1127);
	or gate_anoymous_9_n354 (anoymous_9_n354, anoymous_9_n352, anoymous_9_n351);
	xor gate_anoymous_9_n355 (anoymous_9_n355, anoymous_9_n1127, anoymous_9_n353);
	xor gate_anoymous_9_n348 (anoymous_9_n348, anoymous_9_n1095, anoymous_9_n1111);
	and gate_anoymous_9_n347 (anoymous_9_n347, anoymous_9_n1111, anoymous_9_n1095);
	and gate_anoymous_9_n346 (anoymous_9_n346, anoymous_9_n348, anoymous_9_n1079);
	or gate_anoymous_9_n349 (anoymous_9_n349, anoymous_9_n347, anoymous_9_n346);
	xor gate_anoymous_9_n350 (anoymous_9_n350, anoymous_9_n1079, anoymous_9_n348);
	xor gate_anoymous_9_n343 (anoymous_9_n343, anoymous_9_n1143, anoymous_9_n1159);
	and gate_anoymous_9_n342 (anoymous_9_n342, anoymous_9_n1159, anoymous_9_n1143);
	and gate_anoymous_9_n341 (anoymous_9_n341, anoymous_9_n355, anoymous_9_n343);
	or gate_anoymous_9_n344 (anoymous_9_n344, anoymous_9_n342, anoymous_9_n341);
	xor gate_anoymous_9_n345 (anoymous_9_n345, anoymous_9_n343, anoymous_9_n355);
	xor gate_anoymous_9_n338 (anoymous_9_n338, anoymous_9_n384, anoymous_9_n379);
	and gate_anoymous_9_n337 (anoymous_9_n337, anoymous_9_n379, anoymous_9_n384);
	and gate_anoymous_9_n336 (anoymous_9_n336, anoymous_9_n338, anoymous_9_n350);
	or gate_anoymous_9_n339 (anoymous_9_n339, anoymous_9_n337, anoymous_9_n336);
	xor gate_anoymous_9_n340 (anoymous_9_n340, anoymous_9_n350, anoymous_9_n338);
	xor gate_anoymous_9_n333 (anoymous_9_n333, anoymous_9_n345, anoymous_9_n374);
	and gate_anoymous_9_n332 (anoymous_9_n332, anoymous_9_n374, anoymous_9_n345);
	and gate_anoymous_9_n331 (anoymous_9_n331, anoymous_9_n369, anoymous_9_n333);
	or gate_anoymous_9_n334 (anoymous_9_n334, anoymous_9_n332, anoymous_9_n331);
	xor gate_anoymous_9_n335 (anoymous_9_n335, anoymous_9_n333, anoymous_9_n369);
	xor gate_anoymous_9_n328 (anoymous_9_n328, anoymous_9_n340, anoymous_9_n364);
	and gate_anoymous_9_n327 (anoymous_9_n327, anoymous_9_n364, anoymous_9_n340);
	and gate_anoymous_9_n326 (anoymous_9_n326, anoymous_9_n328, anoymous_9_n335);
	or gate_anoymous_9_n329 (anoymous_9_n329, anoymous_9_n327, anoymous_9_n326);
	xor gate_anoymous_9_n330 (anoymous_9_n330, anoymous_9_n335, anoymous_9_n328);
	not gate_anoymous_9_n325 (anoymous_9_n325, anoymous_9_n324);
	xor gate_anoymous_9_n321 (anoymous_9_n321, anoymous_9_n325, anoymous_9_n1142);
	and gate_anoymous_9_n320 (anoymous_9_n320, anoymous_9_n1142, anoymous_9_n325);
	and gate_anoymous_9_n319 (anoymous_9_n319, anoymous_9_n321, anoymous_9_n1126);
	or gate_anoymous_9_n322 (anoymous_9_n322, anoymous_9_n320, anoymous_9_n319);
	xor gate_anoymous_9_n323 (anoymous_9_n323, anoymous_9_n1126, anoymous_9_n321);
	xor gate_anoymous_9_n316 (anoymous_9_n316, anoymous_9_n1110, anoymous_9_n1094);
	and gate_anoymous_9_n315 (anoymous_9_n315, anoymous_9_n1094, anoymous_9_n1110);
	and gate_anoymous_9_n314 (anoymous_9_n314, anoymous_9_n316, anoymous_9_n1078);
	or gate_anoymous_9_n317 (anoymous_9_n317, anoymous_9_n315, anoymous_9_n314);
	xor gate_anoymous_9_n318 (anoymous_9_n318, anoymous_9_n1078, anoymous_9_n316);
	xor gate_anoymous_9_n311 (anoymous_9_n311, anoymous_9_n354, anoymous_9_n349);
	and gate_anoymous_9_n310 (anoymous_9_n310, anoymous_9_n349, anoymous_9_n354);
	and gate_anoymous_9_n309 (anoymous_9_n309, anoymous_9_n311, anoymous_9_n344);
	or gate_anoymous_9_n312 (anoymous_9_n312, anoymous_9_n310, anoymous_9_n309);
	xor gate_anoymous_9_n313 (anoymous_9_n313, anoymous_9_n344, anoymous_9_n311);
	xor gate_anoymous_9_n306 (anoymous_9_n306, anoymous_9_n323, anoymous_9_n318);
	and gate_anoymous_9_n305 (anoymous_9_n305, anoymous_9_n318, anoymous_9_n323);
	and gate_anoymous_9_n304 (anoymous_9_n304, anoymous_9_n339, anoymous_9_n306);
	or gate_anoymous_9_n307 (anoymous_9_n307, anoymous_9_n305, anoymous_9_n304);
	xor gate_anoymous_9_n308 (anoymous_9_n308, anoymous_9_n306, anoymous_9_n339);
	xor gate_anoymous_9_n301 (anoymous_9_n301, anoymous_9_n313, anoymous_9_n334);
	and gate_anoymous_9_n300 (anoymous_9_n300, anoymous_9_n334, anoymous_9_n313);
	and gate_anoymous_9_n299 (anoymous_9_n299, anoymous_9_n301, anoymous_9_n308);
	or gate_anoymous_9_n302 (anoymous_9_n302, anoymous_9_n300, anoymous_9_n299);
	xor gate_anoymous_9_n303 (anoymous_9_n303, anoymous_9_n308, anoymous_9_n301);
	xor gate_anoymous_9_n296 (anoymous_9_n296, anoymous_9_n324, anoymous_9_n1064);
	and gate_anoymous_9_n295 (anoymous_9_n295, anoymous_9_n1064, anoymous_9_n324);
	and gate_anoymous_9_n294 (anoymous_9_n294, anoymous_9_n296, anoymous_9_n1109);
	or gate_anoymous_9_n297 (anoymous_9_n297, anoymous_9_n295, anoymous_9_n294);
	xor gate_anoymous_9_n298 (anoymous_9_n298, anoymous_9_n1109, anoymous_9_n296);
	xor gate_anoymous_9_n291 (anoymous_9_n291, anoymous_9_n1093, anoymous_9_n1077);
	and gate_anoymous_9_n290 (anoymous_9_n290, anoymous_9_n1077, anoymous_9_n1093);
	and gate_anoymous_9_n289 (anoymous_9_n289, anoymous_9_n291, anoymous_9_n1125);
	or gate_anoymous_9_n292 (anoymous_9_n292, anoymous_9_n290, anoymous_9_n289);
	xor gate_anoymous_9_n293 (anoymous_9_n293, anoymous_9_n1125, anoymous_9_n291);
	xor gate_anoymous_9_n286 (anoymous_9_n286, anoymous_9_n1141, anoymous_9_n298);
	and gate_anoymous_9_n285 (anoymous_9_n285, anoymous_9_n298, anoymous_9_n1141);
	and gate_anoymous_9_n284 (anoymous_9_n284, anoymous_9_n286, anoymous_9_n322);
	or gate_anoymous_9_n287 (anoymous_9_n287, anoymous_9_n285, anoymous_9_n284);
	xor gate_anoymous_9_n288 (anoymous_9_n288, anoymous_9_n322, anoymous_9_n286);
	xor gate_anoymous_9_n281 (anoymous_9_n281, anoymous_9_n317, anoymous_9_n293);
	and gate_anoymous_9_n280 (anoymous_9_n280, anoymous_9_n293, anoymous_9_n317);
	and gate_anoymous_9_n279 (anoymous_9_n279, anoymous_9_n288, anoymous_9_n281);
	or gate_anoymous_9_n282 (anoymous_9_n282, anoymous_9_n280, anoymous_9_n279);
	xor gate_anoymous_9_n283 (anoymous_9_n283, anoymous_9_n281, anoymous_9_n288);
	xor gate_anoymous_9_n276 (anoymous_9_n276, anoymous_9_n312, anoymous_9_n307);
	and gate_anoymous_9_n275 (anoymous_9_n275, anoymous_9_n307, anoymous_9_n312);
	and gate_anoymous_9_n274 (anoymous_9_n274, anoymous_9_n276, anoymous_9_n283);
	or gate_anoymous_9_n277 (anoymous_9_n277, anoymous_9_n275, anoymous_9_n274);
	xor gate_anoymous_9_n278 (anoymous_9_n278, anoymous_9_n283, anoymous_9_n276);
	not gate_anoymous_9_n273 (anoymous_9_n273, anoymous_9_n272);
	xor gate_anoymous_9_n269 (anoymous_9_n269, anoymous_9_n273, anoymous_9_n1124);
	and gate_anoymous_9_n268 (anoymous_9_n268, anoymous_9_n1124, anoymous_9_n273);
	and gate_anoymous_9_n267 (anoymous_9_n267, anoymous_9_n269, anoymous_9_n1108);
	or gate_anoymous_9_n270 (anoymous_9_n270, anoymous_9_n268, anoymous_9_n267);
	xor gate_anoymous_9_n271 (anoymous_9_n271, anoymous_9_n1108, anoymous_9_n269);
	xor gate_anoymous_9_n264 (anoymous_9_n264, anoymous_9_n1092, anoymous_9_n1076);
	and gate_anoymous_9_n263 (anoymous_9_n263, anoymous_9_n1076, anoymous_9_n1092);
	and gate_anoymous_9_n262 (anoymous_9_n262, anoymous_9_n264, anoymous_9_n297);
	or gate_anoymous_9_n265 (anoymous_9_n265, anoymous_9_n263, anoymous_9_n262);
	xor gate_anoymous_9_n266 (anoymous_9_n266, anoymous_9_n297, anoymous_9_n264);
	xor gate_anoymous_9_n259 (anoymous_9_n259, anoymous_9_n292, anoymous_9_n271);
	and gate_anoymous_9_n258 (anoymous_9_n258, anoymous_9_n271, anoymous_9_n292);
	and gate_anoymous_9_n257 (anoymous_9_n257, anoymous_9_n259, anoymous_9_n266);
	or gate_anoymous_9_n260 (anoymous_9_n260, anoymous_9_n258, anoymous_9_n257);
	xor gate_anoymous_9_n261 (anoymous_9_n261, anoymous_9_n266, anoymous_9_n259);
	xor gate_anoymous_9_n254 (anoymous_9_n254, anoymous_9_n287, anoymous_9_n282);
	and gate_anoymous_9_n253 (anoymous_9_n253, anoymous_9_n282, anoymous_9_n287);
	and gate_anoymous_9_n252 (anoymous_9_n252, anoymous_9_n254, anoymous_9_n261);
	or gate_anoymous_9_n255 (anoymous_9_n255, anoymous_9_n253, anoymous_9_n252);
	xor gate_anoymous_9_n256 (anoymous_9_n256, anoymous_9_n261, anoymous_9_n254);
	xor gate_anoymous_9_n249 (anoymous_9_n249, anoymous_9_n272, anoymous_9_n1063);
	and gate_anoymous_9_n248 (anoymous_9_n248, anoymous_9_n1063, anoymous_9_n272);
	and gate_anoymous_9_n247 (anoymous_9_n247, anoymous_9_n249, anoymous_9_n1107);
	or gate_anoymous_9_n250 (anoymous_9_n250, anoymous_9_n248, anoymous_9_n247);
	xor gate_anoymous_9_n251 (anoymous_9_n251, anoymous_9_n1107, anoymous_9_n249);
	xor gate_anoymous_9_n244 (anoymous_9_n244, anoymous_9_n1075, anoymous_9_n1091);
	and gate_anoymous_9_n243 (anoymous_9_n243, anoymous_9_n1091, anoymous_9_n1075);
	and gate_anoymous_9_n242 (anoymous_9_n242, anoymous_9_n244, anoymous_9_n1123);
	or gate_anoymous_9_n245 (anoymous_9_n245, anoymous_9_n243, anoymous_9_n242);
	xor gate_anoymous_9_n246 (anoymous_9_n246, anoymous_9_n1123, anoymous_9_n244);
	xor gate_anoymous_9_n239 (anoymous_9_n239, anoymous_9_n251, anoymous_9_n270);
	and gate_anoymous_9_n238 (anoymous_9_n238, anoymous_9_n270, anoymous_9_n251);
	and gate_anoymous_9_n237 (anoymous_9_n237, anoymous_9_n239, anoymous_9_n265);
	or gate_anoymous_9_n240 (anoymous_9_n240, anoymous_9_n238, anoymous_9_n237);
	xor gate_anoymous_9_n241 (anoymous_9_n241, anoymous_9_n265, anoymous_9_n239);
	xor gate_anoymous_9_n234 (anoymous_9_n234, anoymous_9_n246, anoymous_9_n241);
	and gate_anoymous_9_n233 (anoymous_9_n233, anoymous_9_n241, anoymous_9_n246);
	and gate_anoymous_9_n232 (anoymous_9_n232, anoymous_9_n234, anoymous_9_n260);
	or gate_anoymous_9_n235 (anoymous_9_n235, anoymous_9_n233, anoymous_9_n232);
	xor gate_anoymous_9_n236 (anoymous_9_n236, anoymous_9_n260, anoymous_9_n234);
	not gate_anoymous_9_n231 (anoymous_9_n231, anoymous_9_n230);
	xor gate_anoymous_9_n227 (anoymous_9_n227, anoymous_9_n231, anoymous_9_n1106);
	and gate_anoymous_9_n226 (anoymous_9_n226, anoymous_9_n1106, anoymous_9_n231);
	and gate_anoymous_9_n225 (anoymous_9_n225, anoymous_9_n227, anoymous_9_n1090);
	or gate_anoymous_9_n228 (anoymous_9_n228, anoymous_9_n226, anoymous_9_n225);
	xor gate_anoymous_9_n229 (anoymous_9_n229, anoymous_9_n1090, anoymous_9_n227);
	xor gate_anoymous_9_n222 (anoymous_9_n222, anoymous_9_n1074, anoymous_9_n250);
	and gate_anoymous_9_n221 (anoymous_9_n221, anoymous_9_n250, anoymous_9_n1074);
	and gate_anoymous_9_n220 (anoymous_9_n220, anoymous_9_n245, anoymous_9_n222);
	or gate_anoymous_9_n223 (anoymous_9_n223, anoymous_9_n221, anoymous_9_n220);
	xor gate_anoymous_9_n224 (anoymous_9_n224, anoymous_9_n222, anoymous_9_n245);
	xor gate_anoymous_9_n217 (anoymous_9_n217, anoymous_9_n229, anoymous_9_n224);
	and gate_anoymous_9_n216 (anoymous_9_n216, anoymous_9_n224, anoymous_9_n229);
	and gate_anoymous_9_n215 (anoymous_9_n215, anoymous_9_n217, anoymous_9_n240);
	or gate_anoymous_9_n218 (anoymous_9_n218, anoymous_9_n216, anoymous_9_n215);
	xor gate_anoymous_9_n219 (anoymous_9_n219, anoymous_9_n240, anoymous_9_n217);
	xor gate_anoymous_9_n212 (anoymous_9_n212, anoymous_9_n230, anoymous_9_n1062);
	and gate_anoymous_9_n211 (anoymous_9_n211, anoymous_9_n1062, anoymous_9_n230);
	and gate_anoymous_9_n210 (anoymous_9_n210, anoymous_9_n212, anoymous_9_n1089);
	or gate_anoymous_9_n213 (anoymous_9_n213, anoymous_9_n211, anoymous_9_n210);
	xor gate_anoymous_9_n214 (anoymous_9_n214, anoymous_9_n1089, anoymous_9_n212);
	xor gate_anoymous_9_n207 (anoymous_9_n207, anoymous_9_n1073, anoymous_9_n1105);
	and gate_anoymous_9_n206 (anoymous_9_n206, anoymous_9_n1105, anoymous_9_n1073);
	and gate_anoymous_9_n205 (anoymous_9_n205, anoymous_9_n214, anoymous_9_n207);
	or gate_anoymous_9_n208 (anoymous_9_n208, anoymous_9_n206, anoymous_9_n205);
	xor gate_anoymous_9_n209 (anoymous_9_n209, anoymous_9_n207, anoymous_9_n214);
	xor gate_anoymous_9_n202 (anoymous_9_n202, anoymous_9_n228, anoymous_9_n209);
	and gate_anoymous_9_n201 (anoymous_9_n201, anoymous_9_n209, anoymous_9_n228);
	and gate_anoymous_9_n200 (anoymous_9_n200, anoymous_9_n202, anoymous_9_n223);
	or gate_anoymous_9_n203 (anoymous_9_n203, anoymous_9_n201, anoymous_9_n200);
	xor gate_anoymous_9_n204 (anoymous_9_n204, anoymous_9_n223, anoymous_9_n202);
	not gate_anoymous_9_n199 (anoymous_9_n199, anoymous_9_n198);
	xor gate_anoymous_9_n195 (anoymous_9_n195, anoymous_9_n199, anoymous_9_n1088);
	and gate_anoymous_9_n194 (anoymous_9_n194, anoymous_9_n1088, anoymous_9_n199);
	and gate_anoymous_9_n193 (anoymous_9_n193, anoymous_9_n195, anoymous_9_n1072);
	or gate_anoymous_9_n196 (anoymous_9_n196, anoymous_9_n194, anoymous_9_n193);
	xor gate_anoymous_9_n197 (anoymous_9_n197, anoymous_9_n1072, anoymous_9_n195);
	xor gate_anoymous_9_n190 (anoymous_9_n190, anoymous_9_n213, anoymous_9_n208);
	and gate_anoymous_9_n189 (anoymous_9_n189, anoymous_9_n208, anoymous_9_n213);
	and gate_anoymous_9_n188 (anoymous_9_n188, anoymous_9_n190, anoymous_9_n197);
	or gate_anoymous_9_n191 (anoymous_9_n191, anoymous_9_n189, anoymous_9_n188);
	xor gate_anoymous_9_n192 (anoymous_9_n192, anoymous_9_n197, anoymous_9_n190);
	xor gate_anoymous_9_n185 (anoymous_9_n185, anoymous_9_n198, anoymous_9_n1061);
	and gate_anoymous_9_n184 (anoymous_9_n184, anoymous_9_n1061, anoymous_9_n198);
	and gate_anoymous_9_n183 (anoymous_9_n183, anoymous_9_n185, anoymous_9_n1071);
	or gate_anoymous_9_n186 (anoymous_9_n186, anoymous_9_n184, anoymous_9_n183);
	xor gate_anoymous_9_n187 (anoymous_9_n187, anoymous_9_n1071, anoymous_9_n185);
	xor gate_anoymous_9_n180 (anoymous_9_n180, anoymous_9_n1087, anoymous_9_n187);
	and gate_anoymous_9_n179 (anoymous_9_n179, anoymous_9_n187, anoymous_9_n1087);
	and gate_anoymous_9_n178 (anoymous_9_n178, anoymous_9_n180, anoymous_9_n196);
	or gate_anoymous_9_n181 (anoymous_9_n181, anoymous_9_n179, anoymous_9_n178);
	xor gate_anoymous_9_n182 (anoymous_9_n182, anoymous_9_n196, anoymous_9_n180);
	not gate_anoymous_9_n177 (anoymous_9_n177, anoymous_9_n176);
	xor gate_anoymous_9_n173 (anoymous_9_n173, anoymous_9_n177, anoymous_9_n1070);
	and gate_anoymous_9_n172 (anoymous_9_n172, anoymous_9_n1070, anoymous_9_n177);
	and gate_anoymous_9_n171 (anoymous_9_n171, anoymous_9_n173, anoymous_9_n186);
	or gate_anoymous_9_n174 (anoymous_9_n174, anoymous_9_n172, anoymous_9_n171);
	xor gate_anoymous_9_n175 (anoymous_9_n175, anoymous_9_n186, anoymous_9_n173);
	xor gate_anoymous_9_n169 (anoymous_9_n169, anoymous_9_n1069, anoymous_9_n1060);
	xor gate_anoymous_9_n170 (anoymous_9_n170, anoymous_9_n176, anoymous_9_n169);
	and gate_anoymous_9_n168 (anoymous_9_n168, anoymous_9_n1211, anoymous_9_n1059);
	xor gate_sum_1 (sum_1, anoymous_9_n1059, anoymous_9_n1211);
	xor gate_anoymous_9_n138 (anoymous_9_n138, anoymous_9_n1210, anoymous_9_n1194);
	and gate_anoymous_9_n137 (anoymous_9_n137, anoymous_9_n1194, anoymous_9_n1210);
	and gate_anoymous_9_n136 (anoymous_9_n136, anoymous_9_n138, anoymous_9_n168);
	or gate_anoymous_9_n167 (anoymous_9_n167, anoymous_9_n137, anoymous_9_n136);
	xor gate_sum_2 (sum_2, anoymous_9_n168, anoymous_9_n138);
	xor gate_anoymous_9_n135 (anoymous_9_n135, anoymous_9_n1058, anoymous_9_n754);
	and gate_anoymous_9_n134 (anoymous_9_n134, anoymous_9_n754, anoymous_9_n1058);
	and gate_anoymous_9_n133 (anoymous_9_n133, anoymous_9_n135, anoymous_9_n167);
	or gate_anoymous_9_n166 (anoymous_9_n166, anoymous_9_n134, anoymous_9_n133);
	xor gate_sum_3 (sum_3, anoymous_9_n167, anoymous_9_n135);
	xor gate_anoymous_9_n132 (anoymous_9_n132, anoymous_9_n753, anoymous_9_n752);
	and gate_anoymous_9_n131 (anoymous_9_n131, anoymous_9_n752, anoymous_9_n753);
	and gate_anoymous_9_n130 (anoymous_9_n130, anoymous_9_n132, anoymous_9_n166);
	or gate_anoymous_9_n165 (anoymous_9_n165, anoymous_9_n131, anoymous_9_n130);
	xor gate_sum_4 (sum_4, anoymous_9_n166, anoymous_9_n132);
	xor gate_anoymous_9_n129 (anoymous_9_n129, anoymous_9_n751, anoymous_9_n745);
	and gate_anoymous_9_n128 (anoymous_9_n128, anoymous_9_n745, anoymous_9_n751);
	and gate_anoymous_9_n127 (anoymous_9_n127, anoymous_9_n165, anoymous_9_n129);
	or gate_anoymous_9_n164 (anoymous_9_n164, anoymous_9_n128, anoymous_9_n127);
	xor gate_sum_5 (sum_5, anoymous_9_n129, anoymous_9_n165);
	xor gate_anoymous_9_n126 (anoymous_9_n126, anoymous_9_n740, anoymous_9_n735);
	and gate_anoymous_9_n125 (anoymous_9_n125, anoymous_9_n735, anoymous_9_n740);
	and gate_anoymous_9_n124 (anoymous_9_n124, anoymous_9_n164, anoymous_9_n126);
	or gate_anoymous_9_n163 (anoymous_9_n163, anoymous_9_n125, anoymous_9_n124);
	xor gate_sum_6 (sum_6, anoymous_9_n126, anoymous_9_n164);
	xor gate_anoymous_9_n123 (anoymous_9_n123, anoymous_9_n734, anoymous_9_n723);
	and gate_anoymous_9_n122 (anoymous_9_n122, anoymous_9_n723, anoymous_9_n734);
	and gate_anoymous_9_n121 (anoymous_9_n121, anoymous_9_n163, anoymous_9_n123);
	or gate_anoymous_9_n162 (anoymous_9_n162, anoymous_9_n122, anoymous_9_n121);
	xor gate_sum_7 (sum_7, anoymous_9_n123, anoymous_9_n163);
	xor gate_anoymous_9_n120 (anoymous_9_n120, anoymous_9_n722, anoymous_9_n708);
	and gate_anoymous_9_n119 (anoymous_9_n119, anoymous_9_n708, anoymous_9_n722);
	and gate_anoymous_9_n118 (anoymous_9_n118, anoymous_9_n162, anoymous_9_n120);
	or gate_anoymous_9_n161 (anoymous_9_n161, anoymous_9_n119, anoymous_9_n118);
	xor gate_sum_8 (sum_8, anoymous_9_n120, anoymous_9_n162);
	xor gate_anoymous_9_n117 (anoymous_9_n117, anoymous_9_n707, anoymous_9_n691);
	and gate_anoymous_9_n116 (anoymous_9_n116, anoymous_9_n691, anoymous_9_n707);
	and gate_anoymous_9_n115 (anoymous_9_n115, anoymous_9_n161, anoymous_9_n117);
	or gate_anoymous_9_n160 (anoymous_9_n160, anoymous_9_n116, anoymous_9_n115);
	xor gate_sum_9 (sum_9, anoymous_9_n117, anoymous_9_n161);
	xor gate_anoymous_9_n114 (anoymous_9_n114, anoymous_9_n690, anoymous_9_n671);
	and gate_anoymous_9_n113 (anoymous_9_n113, anoymous_9_n671, anoymous_9_n690);
	and gate_anoymous_9_n112 (anoymous_9_n112, anoymous_9_n160, anoymous_9_n114);
	or gate_anoymous_9_n159 (anoymous_9_n159, anoymous_9_n113, anoymous_9_n112);
	xor gate_sum_10 (sum_10, anoymous_9_n114, anoymous_9_n160);
	xor gate_anoymous_9_n111 (anoymous_9_n111, anoymous_9_n670, anoymous_9_n649);
	and gate_anoymous_9_n110 (anoymous_9_n110, anoymous_9_n649, anoymous_9_n670);
	and gate_anoymous_9_n109 (anoymous_9_n109, anoymous_9_n159, anoymous_9_n111);
	or gate_anoymous_9_n158 (anoymous_9_n158, anoymous_9_n110, anoymous_9_n109);
	xor gate_sum_11 (sum_11, anoymous_9_n111, anoymous_9_n159);
	xor gate_anoymous_9_n108 (anoymous_9_n108, anoymous_9_n648, anoymous_9_n624);
	and gate_anoymous_9_n107 (anoymous_9_n107, anoymous_9_n624, anoymous_9_n648);
	and gate_anoymous_9_n106 (anoymous_9_n106, anoymous_9_n158, anoymous_9_n108);
	or gate_anoymous_9_n157 (anoymous_9_n157, anoymous_9_n107, anoymous_9_n106);
	xor gate_sum_12 (sum_12, anoymous_9_n108, anoymous_9_n158);
	xor gate_anoymous_9_n105 (anoymous_9_n105, anoymous_9_n623, anoymous_9_n597);
	and gate_anoymous_9_n104 (anoymous_9_n104, anoymous_9_n597, anoymous_9_n623);
	and gate_anoymous_9_n103 (anoymous_9_n103, anoymous_9_n157, anoymous_9_n105);
	or gate_anoymous_9_n156 (anoymous_9_n156, anoymous_9_n104, anoymous_9_n103);
	xor gate_sum_13 (sum_13, anoymous_9_n105, anoymous_9_n157);
	xor gate_anoymous_9_n102 (anoymous_9_n102, anoymous_9_n596, anoymous_9_n567);
	and gate_anoymous_9_n101 (anoymous_9_n101, anoymous_9_n567, anoymous_9_n596);
	and gate_anoymous_9_n100 (anoymous_9_n100, anoymous_9_n156, anoymous_9_n102);
	or gate_anoymous_9_n155 (anoymous_9_n155, anoymous_9_n101, anoymous_9_n100);
	xor gate_sum_14 (sum_14, anoymous_9_n102, anoymous_9_n156);
	xor gate_anoymous_9_n99 (anoymous_9_n99, anoymous_9_n566, anoymous_9_n535);
	and gate_anoymous_9_n98 (anoymous_9_n98, anoymous_9_n535, anoymous_9_n566);
	and gate_anoymous_9_n97 (anoymous_9_n97, anoymous_9_n155, anoymous_9_n99);
	or gate_anoymous_9_n154 (anoymous_9_n154, anoymous_9_n98, anoymous_9_n97);
	xor gate_sum_15 (sum_15, anoymous_9_n99, anoymous_9_n155);
	xor gate_anoymous_9_n96 (anoymous_9_n96, anoymous_9_n534, anoymous_9_n500);
	and gate_anoymous_9_n95 (anoymous_9_n95, anoymous_9_n500, anoymous_9_n534);
	and gate_anoymous_9_n94 (anoymous_9_n94, anoymous_9_n154, anoymous_9_n96);
	or gate_anoymous_9_n153 (anoymous_9_n153, anoymous_9_n95, anoymous_9_n94);
	xor gate_sum_16 (sum_16, anoymous_9_n96, anoymous_9_n154);
	xor gate_anoymous_9_n93 (anoymous_9_n93, anoymous_9_n499, anoymous_9_n464);
	and gate_anoymous_9_n92 (anoymous_9_n92, anoymous_9_n464, anoymous_9_n499);
	and gate_anoymous_9_n91 (anoymous_9_n91, anoymous_9_n153, anoymous_9_n93);
	or gate_anoymous_9_n152 (anoymous_9_n152, anoymous_9_n92, anoymous_9_n91);
	xor gate_sum_17 (sum_17, anoymous_9_n93, anoymous_9_n153);
	xor gate_anoymous_9_n90 (anoymous_9_n90, anoymous_9_n463, anoymous_9_n427);
	and gate_anoymous_9_n89 (anoymous_9_n89, anoymous_9_n427, anoymous_9_n463);
	and gate_anoymous_9_n88 (anoymous_9_n88, anoymous_9_n152, anoymous_9_n90);
	or gate_anoymous_9_n151 (anoymous_9_n151, anoymous_9_n89, anoymous_9_n88);
	xor gate_sum_18 (sum_18, anoymous_9_n90, anoymous_9_n152);
	xor gate_anoymous_9_n87 (anoymous_9_n87, anoymous_9_n426, anoymous_9_n392);
	and gate_anoymous_9_n86 (anoymous_9_n86, anoymous_9_n392, anoymous_9_n426);
	and gate_anoymous_9_n85 (anoymous_9_n85, anoymous_9_n151, anoymous_9_n87);
	or gate_anoymous_9_n150 (anoymous_9_n150, anoymous_9_n86, anoymous_9_n85);
	xor gate_sum_19 (sum_19, anoymous_9_n87, anoymous_9_n151);
	xor gate_anoymous_9_n84 (anoymous_9_n84, anoymous_9_n391, anoymous_9_n360);
	and gate_anoymous_9_n83 (anoymous_9_n83, anoymous_9_n360, anoymous_9_n391);
	and gate_anoymous_9_n82 (anoymous_9_n82, anoymous_9_n150, anoymous_9_n84);
	or gate_anoymous_9_n149 (anoymous_9_n149, anoymous_9_n83, anoymous_9_n82);
	xor gate_sum_20 (sum_20, anoymous_9_n84, anoymous_9_n150);
	xor gate_anoymous_9_n81 (anoymous_9_n81, anoymous_9_n359, anoymous_9_n330);
	and gate_anoymous_9_n80 (anoymous_9_n80, anoymous_9_n330, anoymous_9_n359);
	and gate_anoymous_9_n79 (anoymous_9_n79, anoymous_9_n149, anoymous_9_n81);
	or gate_anoymous_9_n148 (anoymous_9_n148, anoymous_9_n80, anoymous_9_n79);
	xor gate_sum_21 (sum_21, anoymous_9_n81, anoymous_9_n149);
	xor gate_anoymous_9_n78 (anoymous_9_n78, anoymous_9_n329, anoymous_9_n303);
	and gate_anoymous_9_n77 (anoymous_9_n77, anoymous_9_n303, anoymous_9_n329);
	and gate_anoymous_9_n76 (anoymous_9_n76, anoymous_9_n148, anoymous_9_n78);
	or gate_anoymous_9_n147 (anoymous_9_n147, anoymous_9_n77, anoymous_9_n76);
	xor gate_sum_22 (sum_22, anoymous_9_n78, anoymous_9_n148);
	xor gate_anoymous_9_n75 (anoymous_9_n75, anoymous_9_n302, anoymous_9_n278);
	and gate_anoymous_9_n74 (anoymous_9_n74, anoymous_9_n278, anoymous_9_n302);
	and gate_anoymous_9_n73 (anoymous_9_n73, anoymous_9_n147, anoymous_9_n75);
	or gate_anoymous_9_n146 (anoymous_9_n146, anoymous_9_n74, anoymous_9_n73);
	xor gate_sum_23 (sum_23, anoymous_9_n75, anoymous_9_n147);
	xor gate_anoymous_9_n72 (anoymous_9_n72, anoymous_9_n277, anoymous_9_n256);
	and gate_anoymous_9_n71 (anoymous_9_n71, anoymous_9_n256, anoymous_9_n277);
	and gate_anoymous_9_n70 (anoymous_9_n70, anoymous_9_n146, anoymous_9_n72);
	or gate_anoymous_9_n145 (anoymous_9_n145, anoymous_9_n71, anoymous_9_n70);
	xor gate_sum_24 (sum_24, anoymous_9_n72, anoymous_9_n146);
	xor gate_anoymous_9_n69 (anoymous_9_n69, anoymous_9_n255, anoymous_9_n236);
	and gate_anoymous_9_n68 (anoymous_9_n68, anoymous_9_n236, anoymous_9_n255);
	and gate_anoymous_9_n67 (anoymous_9_n67, anoymous_9_n145, anoymous_9_n69);
	or gate_anoymous_9_n144 (anoymous_9_n144, anoymous_9_n68, anoymous_9_n67);
	xor gate_sum_25 (sum_25, anoymous_9_n69, anoymous_9_n145);
	xor gate_anoymous_9_n66 (anoymous_9_n66, anoymous_9_n219, anoymous_9_n235);
	and gate_anoymous_9_n65 (anoymous_9_n65, anoymous_9_n235, anoymous_9_n219);
	and gate_anoymous_9_n64 (anoymous_9_n64, anoymous_9_n144, anoymous_9_n66);
	or gate_anoymous_9_n143 (anoymous_9_n143, anoymous_9_n65, anoymous_9_n64);
	xor gate_sum_26 (sum_26, anoymous_9_n66, anoymous_9_n144);
	xor gate_anoymous_9_n63 (anoymous_9_n63, anoymous_9_n204, anoymous_9_n218);
	and gate_anoymous_9_n62 (anoymous_9_n62, anoymous_9_n218, anoymous_9_n204);
	and gate_anoymous_9_n61 (anoymous_9_n61, anoymous_9_n143, anoymous_9_n63);
	or gate_anoymous_9_n142 (anoymous_9_n142, anoymous_9_n62, anoymous_9_n61);
	xor gate_sum_27 (sum_27, anoymous_9_n63, anoymous_9_n143);
	xor gate_anoymous_9_n60 (anoymous_9_n60, anoymous_9_n203, anoymous_9_n192);
	and gate_anoymous_9_n59 (anoymous_9_n59, anoymous_9_n192, anoymous_9_n203);
	and gate_anoymous_9_n58 (anoymous_9_n58, anoymous_9_n142, anoymous_9_n60);
	or gate_anoymous_9_n141 (anoymous_9_n141, anoymous_9_n59, anoymous_9_n58);
	xor gate_sum_28 (sum_28, anoymous_9_n60, anoymous_9_n142);
	xor gate_anoymous_9_n57 (anoymous_9_n57, anoymous_9_n182, anoymous_9_n191);
	and gate_anoymous_9_n56 (anoymous_9_n56, anoymous_9_n191, anoymous_9_n182);
	and gate_anoymous_9_n55 (anoymous_9_n55, anoymous_9_n141, anoymous_9_n57);
	or gate_anoymous_9_n140 (anoymous_9_n140, anoymous_9_n56, anoymous_9_n55);
	xor gate_sum_29 (sum_29, anoymous_9_n57, anoymous_9_n141);
	xor gate_anoymous_9_n54 (anoymous_9_n54, anoymous_9_n175, anoymous_9_n181);
	and gate_anoymous_9_n53 (anoymous_9_n53, anoymous_9_n181, anoymous_9_n175);
	and gate_anoymous_9_n52 (anoymous_9_n52, anoymous_9_n140, anoymous_9_n54);
	or gate_anoymous_9_n139 (anoymous_9_n139, anoymous_9_n53, anoymous_9_n52);
	xor gate_sum_30 (sum_30, anoymous_9_n54, anoymous_9_n140);
	xor gate_anoymous_9_n51 (anoymous_9_n51, anoymous_9_n170, anoymous_9_n174);
	xor gate_sum_31 (sum_31, anoymous_9_n51, anoymous_9_n139);
	buf gate_anoymous_9_n49 (anoymous_9_n49, b_0);
	buf gate_anoymous_9_n48 (anoymous_9_n48, anoymous_9_n1387);
	buf gate_anoymous_9_n47 (anoymous_9_n47, anoymous_9_n1387);
	buf gate_anoymous_9_n46 (anoymous_9_n46, anoymous_9_n1396);
	buf gate_anoymous_9_n45 (anoymous_9_n45, anoymous_9_n1396);
	buf gate_anoymous_9_n43 (anoymous_9_n43, a_15);
	buf gate_anoymous_9_n42 (anoymous_9_n42, anoymous_9_n1388);
	buf gate_anoymous_9_n41 (anoymous_9_n41, anoymous_9_n1388);
	buf gate_anoymous_9_n40 (anoymous_9_n40, anoymous_9_n1397);
	buf gate_anoymous_9_n39 (anoymous_9_n39, anoymous_9_n1397);
	buf gate_anoymous_9_n37 (anoymous_9_n37, a_13);
	buf gate_anoymous_9_n36 (anoymous_9_n36, anoymous_9_n1389);
	buf gate_anoymous_9_n35 (anoymous_9_n35, anoymous_9_n1389);
	buf gate_anoymous_9_n34 (anoymous_9_n34, anoymous_9_n1398);
	buf gate_anoymous_9_n33 (anoymous_9_n33, anoymous_9_n1398);
	buf gate_anoymous_9_n31 (anoymous_9_n31, a_11);
	buf gate_anoymous_9_n30 (anoymous_9_n30, anoymous_9_n1390);
	buf gate_anoymous_9_n29 (anoymous_9_n29, anoymous_9_n1390);
	buf gate_anoymous_9_n28 (anoymous_9_n28, anoymous_9_n1399);
	buf gate_anoymous_9_n27 (anoymous_9_n27, anoymous_9_n1399);
	buf gate_anoymous_9_n25 (anoymous_9_n25, a_9);
	buf gate_anoymous_9_n24 (anoymous_9_n24, anoymous_9_n1391);
	buf gate_anoymous_9_n23 (anoymous_9_n23, anoymous_9_n1391);
	buf gate_anoymous_9_n22 (anoymous_9_n22, anoymous_9_n1400);
	buf gate_anoymous_9_n21 (anoymous_9_n21, anoymous_9_n1400);
	buf gate_anoymous_9_n19 (anoymous_9_n19, a_7);
	buf gate_anoymous_9_n18 (anoymous_9_n18, anoymous_9_n1392);
	buf gate_anoymous_9_n17 (anoymous_9_n17, anoymous_9_n1392);
	buf gate_anoymous_9_n16 (anoymous_9_n16, anoymous_9_n1401);
	buf gate_anoymous_9_n15 (anoymous_9_n15, anoymous_9_n1401);
	buf gate_anoymous_9_n13 (anoymous_9_n13, a_5);
	buf gate_anoymous_9_n12 (anoymous_9_n12, anoymous_9_n1393);
	buf gate_anoymous_9_n11 (anoymous_9_n11, anoymous_9_n1393);
	buf gate_anoymous_9_n10 (anoymous_9_n10, anoymous_9_n1402);
	buf gate_anoymous_9_n9 (anoymous_9_n9, anoymous_9_n1402);
	buf gate_anoymous_9_n7 (anoymous_9_n7, a_3);
	buf gate_anoymous_9_n6 (anoymous_9_n6, anoymous_9_n1394);
	buf gate_anoymous_9_n5 (anoymous_9_n5, anoymous_9_n1394);
	buf gate_anoymous_9_n4 (anoymous_9_n4, anoymous_9_n1403);
	buf gate_anoymous_9_n3 (anoymous_9_n3, anoymous_9_n1403);
	buf gate_anoymous_9_n1 (anoymous_9_n1, a_1);
endmodule

