
module multiplier_16_bit (a_0, a_1, a_2, a_3, a_4, a_5, a_6, a_7, a_8, a_9, a_10, a_11, a_12, a_13, a_14, a_15, 
   b_0, b_1, b_2, b_3, b_4, b_5, b_6, b_7, b_8, b_9, b_10, b_11, b_12, b_13, b_14, b_15,
   sum_0, sum_1, sum_2, sum_3, sum_4, sum_5, sum_6, sum_7, sum_8, sum_9, sum_10, sum_11, 
   sum_12, sum_13, sum_14, sum_15, sum_16, sum_17, sum_18, sum_19, sum_20, sum_21, sum_22, 
   sum_23, sum_24, sum_25, sum_26, sum_27, sum_28, sum_29, sum_30, sum_31);

  input a_0;
  input a_1;
  input a_2;
  input a_3;
  input a_4;
  input a_5;
  input a_6;
  input a_7;
  input a_8;
  input a_9;
  input a_10;
  input a_11;
  input a_12;
  input a_13;
  input a_14;
  input a_15;

  input b_0;
  input b_1;
  input b_2;
  input b_3;
  input b_4;
  input b_5;
  input b_6;
  input b_7;
  input b_8;
  input b_9;
  input b_10;
  input b_11;
  input b_12;
  input b_13;
  input b_14;
  input b_15;


  output sum_0;
  output sum_1;
  output sum_2;
  output sum_3;
  output sum_4;
  output sum_5;
  output sum_6;
  output sum_7;
  output sum_8;
  output sum_9;
  output sum_10;
  output sum_11;
  output sum_12;
  output sum_13;
  output sum_14;
  output sum_15;
  output sum_16;
output sum_17;
output sum_18;
output sum_19;
output sum_20;
output sum_21;
output sum_22;
output sum_23;
output sum_24;
output sum_25;
output sum_26;
output sum_27;
output sum_28;
output sum_29;
output sum_30;
output sum_31;
  

	not gate_mult_9_n1403 (mult_9_n1403, a_0);
	xor gate_mult_9_n1386 (mult_9_n1386, a_1, a_0);
	nand gate_mult_9_n1394 (mult_9_n1394, mult_9_n1403, mult_9_n1386);
	xnor gate_mult_9_n1402 (mult_9_n1402, a_1, a_2);
	xor gate_mult_9_n1385 (mult_9_n1385, a_3, a_2);
	nand gate_mult_9_n1393 (mult_9_n1393, mult_9_n1385, mult_9_n1402);
	xnor gate_mult_9_n1401 (mult_9_n1401, a_3, a_4);
	xor gate_mult_9_n1384 (mult_9_n1384, a_5, a_4);
	nand gate_mult_9_n1392 (mult_9_n1392, mult_9_n1384, mult_9_n1401);
	xnor gate_mult_9_n1400 (mult_9_n1400, a_5, a_6);
	xor gate_mult_9_n1383 (mult_9_n1383, a_7, a_6);
	nand gate_mult_9_n1391 (mult_9_n1391, mult_9_n1383, mult_9_n1400);
	xnor gate_mult_9_n1399 (mult_9_n1399, a_7, a_8);
	xor gate_mult_9_n1382 (mult_9_n1382, a_9, a_8);
	nand gate_mult_9_n1390 (mult_9_n1390, mult_9_n1382, mult_9_n1399);
	xnor gate_mult_9_n1398 (mult_9_n1398, a_9, a_10);
	xor gate_mult_9_n1381 (mult_9_n1381, a_11, a_10);
	nand gate_mult_9_n1389 (mult_9_n1389, mult_9_n1381, mult_9_n1398);
	xnor gate_mult_9_n1397 (mult_9_n1397, a_11, a_12);
	xor gate_mult_9_n1380 (mult_9_n1380, a_13, a_12);
	nand gate_mult_9_n1388 (mult_9_n1388, mult_9_n1380, mult_9_n1397);
	xnor gate_mult_9_n1396 (mult_9_n1396, a_13, a_14);
	xor gate_mult_9_n1379 (mult_9_n1379, a_15, a_14);
	nand gate_mult_9_n1387 (mult_9_n1387, mult_9_n1379, mult_9_n1396);
	not gate_mult_9_n1420 (mult_9_n1420, a_15);
	not gate_mult_9_n1411 (mult_9_n1411, mult_9_n1);
	not gate_mult_9_n1410 (mult_9_n1410, mult_9_n7);
	not gate_mult_9_n1409 (mult_9_n1409, mult_9_n13);
	not gate_mult_9_n1408 (mult_9_n1408, mult_9_n19);
	not gate_mult_9_n1407 (mult_9_n1407, mult_9_n25);
	not gate_mult_9_n1406 (mult_9_n1406, mult_9_n31);
	not gate_mult_9_n1405 (mult_9_n1405, mult_9_n37);
	not gate_mult_9_n1404 (mult_9_n1404, mult_9_n43);
	buf gate_mult_9_n1395 (mult_9_n1395, mult_9_n1420);
	buf gate_mult_9_n1377 (mult_9_n1377, b_1);
	buf gate_mult_9_n1376 (mult_9_n1376, b_2);
	buf gate_mult_9_n1375 (mult_9_n1375, b_3);
	buf gate_mult_9_n1374 (mult_9_n1374, b_4);
	buf gate_mult_9_n1373 (mult_9_n1373, b_5);
	buf gate_mult_9_n1372 (mult_9_n1372, b_6);
	buf gate_mult_9_n1371 (mult_9_n1371, b_7);
	buf gate_mult_9_n1370 (mult_9_n1370, b_8);
	buf gate_mult_9_n1369 (mult_9_n1369, b_9);
	buf gate_mult_9_n1368 (mult_9_n1368, b_10);
	buf gate_mult_9_n1367 (mult_9_n1367, b_11);
	buf gate_mult_9_n1366 (mult_9_n1366, b_12);
	buf gate_mult_9_n1365 (mult_9_n1365, b_13);
	buf gate_mult_9_n1364 (mult_9_n1364, b_14);
	buf gate_mult_9_n1363 (mult_9_n1363, b_15);
	or gate_mult_9_n1362 (mult_9_n1362, mult_9_n49, mult_9_n1411);
	xnor gate_mult_9_n1361 (mult_9_n1361, mult_9_n49, mult_9_n1);
	xnor gate_mult_9_n1360 (mult_9_n1360, mult_9_n1377, mult_9_n1);
	xnor gate_mult_9_n1359 (mult_9_n1359, mult_9_n1376, mult_9_n1);
	xnor gate_mult_9_n1358 (mult_9_n1358, mult_9_n1375, mult_9_n1);
	xnor gate_mult_9_n1357 (mult_9_n1357, mult_9_n1374, mult_9_n1);
	xnor gate_mult_9_n1356 (mult_9_n1356, mult_9_n1373, mult_9_n1);
	xnor gate_mult_9_n1355 (mult_9_n1355, mult_9_n1372, mult_9_n1);
	xnor gate_mult_9_n1354 (mult_9_n1354, mult_9_n1371, mult_9_n1);
	xnor gate_mult_9_n1353 (mult_9_n1353, mult_9_n1370, mult_9_n1);
	xnor gate_mult_9_n1352 (mult_9_n1352, mult_9_n1369, mult_9_n1);
	xnor gate_mult_9_n1351 (mult_9_n1351, mult_9_n1368, mult_9_n1);
	xnor gate_mult_9_n1350 (mult_9_n1350, mult_9_n1367, mult_9_n1);
	xnor gate_mult_9_n1349 (mult_9_n1349, mult_9_n1366, mult_9_n1);
	xnor gate_mult_9_n1348 (mult_9_n1348, mult_9_n1365, mult_9_n1);
	xnor gate_mult_9_n1347 (mult_9_n1347, mult_9_n1364, mult_9_n1);
	xnor gate_mult_9_n1346 (mult_9_n1346, mult_9_n1363, mult_9_n1);
	not gate_mult_9_n1050 (mult_9_n1050, mult_9_n3);
	and gate_sum_0 (sum_0, mult_9_n49, mult_9_n1050);
	or gate_mult_9_n1049 (mult_9_n1049, mult_9_n5, mult_9_n1361);
	or gate_mult_9_n1048 (mult_9_n1048, mult_9_n1360, mult_9_n3);
	nand gate_mult_9_n1211 (mult_9_n1211, mult_9_n1049, mult_9_n1048);
	or gate_mult_9_n1047 (mult_9_n1047, mult_9_n5, mult_9_n1360);
	or gate_mult_9_n1046 (mult_9_n1046, mult_9_n1359, mult_9_n3);
	nand gate_mult_9_n1210 (mult_9_n1210, mult_9_n1047, mult_9_n1046);
	or gate_mult_9_n1045 (mult_9_n1045, mult_9_n5, mult_9_n1359);
	or gate_mult_9_n1044 (mult_9_n1044, mult_9_n1358, mult_9_n3);
	nand gate_mult_9_n1209 (mult_9_n1209, mult_9_n1045, mult_9_n1044);
	or gate_mult_9_n1043 (mult_9_n1043, mult_9_n5, mult_9_n1358);
	or gate_mult_9_n1042 (mult_9_n1042, mult_9_n1357, mult_9_n3);
	nand gate_mult_9_n1208 (mult_9_n1208, mult_9_n1043, mult_9_n1042);
	or gate_mult_9_n1041 (mult_9_n1041, mult_9_n5, mult_9_n1357);
	or gate_mult_9_n1040 (mult_9_n1040, mult_9_n1356, mult_9_n3);
	nand gate_mult_9_n1207 (mult_9_n1207, mult_9_n1041, mult_9_n1040);
	or gate_mult_9_n1039 (mult_9_n1039, mult_9_n5, mult_9_n1356);
	or gate_mult_9_n1038 (mult_9_n1038, mult_9_n1355, mult_9_n3);
	nand gate_mult_9_n1206 (mult_9_n1206, mult_9_n1039, mult_9_n1038);
	or gate_mult_9_n1037 (mult_9_n1037, mult_9_n5, mult_9_n1355);
	or gate_mult_9_n1036 (mult_9_n1036, mult_9_n1354, mult_9_n3);
	nand gate_mult_9_n1205 (mult_9_n1205, mult_9_n1037, mult_9_n1036);
	or gate_mult_9_n1035 (mult_9_n1035, mult_9_n5, mult_9_n1354);
	or gate_mult_9_n1034 (mult_9_n1034, mult_9_n1353, mult_9_n3);
	nand gate_mult_9_n1204 (mult_9_n1204, mult_9_n1035, mult_9_n1034);
	or gate_mult_9_n1033 (mult_9_n1033, mult_9_n5, mult_9_n1353);
	or gate_mult_9_n1032 (mult_9_n1032, mult_9_n1352, mult_9_n4);
	nand gate_mult_9_n1203 (mult_9_n1203, mult_9_n1033, mult_9_n1032);
	or gate_mult_9_n1031 (mult_9_n1031, mult_9_n6, mult_9_n1352);
	or gate_mult_9_n1030 (mult_9_n1030, mult_9_n1351, mult_9_n4);
	nand gate_mult_9_n1202 (mult_9_n1202, mult_9_n1031, mult_9_n1030);
	or gate_mult_9_n1029 (mult_9_n1029, mult_9_n6, mult_9_n1351);
	or gate_mult_9_n1028 (mult_9_n1028, mult_9_n1350, mult_9_n4);
	nand gate_mult_9_n1201 (mult_9_n1201, mult_9_n1029, mult_9_n1028);
	or gate_mult_9_n1027 (mult_9_n1027, mult_9_n6, mult_9_n1350);
	or gate_mult_9_n1026 (mult_9_n1026, mult_9_n1349, mult_9_n4);
	nand gate_mult_9_n1200 (mult_9_n1200, mult_9_n1027, mult_9_n1026);
	or gate_mult_9_n1025 (mult_9_n1025, mult_9_n6, mult_9_n1349);
	or gate_mult_9_n1024 (mult_9_n1024, mult_9_n1348, mult_9_n4);
	nand gate_mult_9_n1199 (mult_9_n1199, mult_9_n1025, mult_9_n1024);
	or gate_mult_9_n1023 (mult_9_n1023, mult_9_n6, mult_9_n1348);
	or gate_mult_9_n1022 (mult_9_n1022, mult_9_n1347, mult_9_n4);
	nand gate_mult_9_n1198 (mult_9_n1198, mult_9_n1023, mult_9_n1022);
	or gate_mult_9_n1021 (mult_9_n1021, mult_9_n6, mult_9_n1347);
	or gate_mult_9_n1020 (mult_9_n1020, mult_9_n1346, mult_9_n4);
	nand gate_mult_9_n1197 (mult_9_n1197, mult_9_n1021, mult_9_n1020);
	or gate_mult_9_n1019 (mult_9_n1019, mult_9_n6, mult_9_n1346);
	or gate_mult_9_n1018 (mult_9_n1018, mult_9_n1411, mult_9_n4);
	nand gate_mult_9_n1196 (mult_9_n1196, mult_9_n1019, mult_9_n1018);
	and gate_mult_9_n1017 (mult_9_n1017, mult_9_n6, mult_9_n4);
	or gate_mult_9_n1195 (mult_9_n1195, mult_9_n1411, mult_9_n1017);
	or gate_mult_9_n1016 (mult_9_n1016, mult_9_n1362, mult_9_n4);
	or gate_mult_9_n1015 (mult_9_n1015, mult_9_n6, mult_9_n1411);
	nand gate_mult_9_n1059 (mult_9_n1059, mult_9_n1016, mult_9_n1015);
	or gate_mult_9_n1345 (mult_9_n1345, mult_9_n49, mult_9_n1410);
	xnor gate_mult_9_n1344 (mult_9_n1344, mult_9_n49, mult_9_n7);
	xnor gate_mult_9_n1343 (mult_9_n1343, mult_9_n1377, mult_9_n7);
	xnor gate_mult_9_n1342 (mult_9_n1342, mult_9_n1376, mult_9_n7);
	xnor gate_mult_9_n1341 (mult_9_n1341, mult_9_n1375, mult_9_n7);
	xnor gate_mult_9_n1340 (mult_9_n1340, mult_9_n1374, mult_9_n7);
	xnor gate_mult_9_n1339 (mult_9_n1339, mult_9_n1373, mult_9_n7);
	xnor gate_mult_9_n1338 (mult_9_n1338, mult_9_n1372, mult_9_n7);
	xnor gate_mult_9_n1337 (mult_9_n1337, mult_9_n1371, mult_9_n7);
	xnor gate_mult_9_n1336 (mult_9_n1336, mult_9_n1370, mult_9_n7);
	xnor gate_mult_9_n1335 (mult_9_n1335, mult_9_n1369, mult_9_n7);
	xnor gate_mult_9_n1334 (mult_9_n1334, mult_9_n1368, mult_9_n7);
	xnor gate_mult_9_n1333 (mult_9_n1333, mult_9_n1367, mult_9_n7);
	xnor gate_mult_9_n1332 (mult_9_n1332, mult_9_n1366, mult_9_n7);
	xnor gate_mult_9_n1331 (mult_9_n1331, mult_9_n1365, mult_9_n7);
	xnor gate_mult_9_n1330 (mult_9_n1330, mult_9_n1364, mult_9_n7);
	xnor gate_mult_9_n1329 (mult_9_n1329, mult_9_n1363, mult_9_n7);
	not gate_mult_9_n1013 (mult_9_n1013, mult_9_n9);
	and gate_mult_9_n1194 (mult_9_n1194, mult_9_n49, mult_9_n1013);
	or gate_mult_9_n1012 (mult_9_n1012, mult_9_n11, mult_9_n1344);
	or gate_mult_9_n1011 (mult_9_n1011, mult_9_n9, mult_9_n1343);
	nand gate_mult_9_n1193 (mult_9_n1193, mult_9_n1012, mult_9_n1011);
	or gate_mult_9_n1010 (mult_9_n1010, mult_9_n11, mult_9_n1343);
	or gate_mult_9_n1009 (mult_9_n1009, mult_9_n9, mult_9_n1342);
	nand gate_mult_9_n1192 (mult_9_n1192, mult_9_n1010, mult_9_n1009);
	or gate_mult_9_n1008 (mult_9_n1008, mult_9_n11, mult_9_n1342);
	or gate_mult_9_n1007 (mult_9_n1007, mult_9_n9, mult_9_n1341);
	nand gate_mult_9_n1191 (mult_9_n1191, mult_9_n1008, mult_9_n1007);
	or gate_mult_9_n1006 (mult_9_n1006, mult_9_n11, mult_9_n1341);
	or gate_mult_9_n1005 (mult_9_n1005, mult_9_n9, mult_9_n1340);
	nand gate_mult_9_n1190 (mult_9_n1190, mult_9_n1006, mult_9_n1005);
	or gate_mult_9_n1004 (mult_9_n1004, mult_9_n11, mult_9_n1340);
	or gate_mult_9_n1003 (mult_9_n1003, mult_9_n9, mult_9_n1339);
	nand gate_mult_9_n1189 (mult_9_n1189, mult_9_n1004, mult_9_n1003);
	or gate_mult_9_n1002 (mult_9_n1002, mult_9_n11, mult_9_n1339);
	or gate_mult_9_n1001 (mult_9_n1001, mult_9_n9, mult_9_n1338);
	nand gate_mult_9_n1188 (mult_9_n1188, mult_9_n1002, mult_9_n1001);
	or gate_mult_9_n1000 (mult_9_n1000, mult_9_n11, mult_9_n1338);
	or gate_mult_9_n999 (mult_9_n999, mult_9_n9, mult_9_n1337);
	nand gate_mult_9_n1187 (mult_9_n1187, mult_9_n1000, mult_9_n999);
	or gate_mult_9_n998 (mult_9_n998, mult_9_n11, mult_9_n1337);
	or gate_mult_9_n997 (mult_9_n997, mult_9_n9, mult_9_n1336);
	nand gate_mult_9_n1186 (mult_9_n1186, mult_9_n998, mult_9_n997);
	or gate_mult_9_n996 (mult_9_n996, mult_9_n11, mult_9_n1336);
	or gate_mult_9_n995 (mult_9_n995, mult_9_n10, mult_9_n1335);
	nand gate_mult_9_n1185 (mult_9_n1185, mult_9_n996, mult_9_n995);
	or gate_mult_9_n994 (mult_9_n994, mult_9_n12, mult_9_n1335);
	or gate_mult_9_n993 (mult_9_n993, mult_9_n10, mult_9_n1334);
	nand gate_mult_9_n1184 (mult_9_n1184, mult_9_n994, mult_9_n993);
	or gate_mult_9_n992 (mult_9_n992, mult_9_n12, mult_9_n1334);
	or gate_mult_9_n991 (mult_9_n991, mult_9_n10, mult_9_n1333);
	nand gate_mult_9_n1183 (mult_9_n1183, mult_9_n992, mult_9_n991);
	or gate_mult_9_n990 (mult_9_n990, mult_9_n12, mult_9_n1333);
	or gate_mult_9_n989 (mult_9_n989, mult_9_n10, mult_9_n1332);
	nand gate_mult_9_n1182 (mult_9_n1182, mult_9_n990, mult_9_n989);
	or gate_mult_9_n988 (mult_9_n988, mult_9_n12, mult_9_n1332);
	or gate_mult_9_n987 (mult_9_n987, mult_9_n10, mult_9_n1331);
	nand gate_mult_9_n1181 (mult_9_n1181, mult_9_n988, mult_9_n987);
	or gate_mult_9_n986 (mult_9_n986, mult_9_n12, mult_9_n1331);
	or gate_mult_9_n985 (mult_9_n985, mult_9_n10, mult_9_n1330);
	nand gate_mult_9_n1180 (mult_9_n1180, mult_9_n986, mult_9_n985);
	or gate_mult_9_n984 (mult_9_n984, mult_9_n12, mult_9_n1330);
	or gate_mult_9_n983 (mult_9_n983, mult_9_n10, mult_9_n1329);
	nand gate_mult_9_n1179 (mult_9_n1179, mult_9_n984, mult_9_n983);
	or gate_mult_9_n982 (mult_9_n982, mult_9_n12, mult_9_n1329);
	or gate_mult_9_n981 (mult_9_n981, mult_9_n10, mult_9_n1410);
	nand gate_mult_9_n1178 (mult_9_n1178, mult_9_n982, mult_9_n981);
	and gate_mult_9_n980 (mult_9_n980, mult_9_n12, mult_9_n10);
	or gate_mult_9_n1177 (mult_9_n1177, mult_9_n1410, mult_9_n980);
	or gate_mult_9_n979 (mult_9_n979, mult_9_n10, mult_9_n1345);
	or gate_mult_9_n978 (mult_9_n978, mult_9_n12, mult_9_n1410);
	nand gate_mult_9_n1058 (mult_9_n1058, mult_9_n979, mult_9_n978);
	or gate_mult_9_n1328 (mult_9_n1328, mult_9_n49, mult_9_n1409);
	xnor gate_mult_9_n1327 (mult_9_n1327, mult_9_n49, mult_9_n13);
	xnor gate_mult_9_n1326 (mult_9_n1326, mult_9_n1377, mult_9_n13);
	xnor gate_mult_9_n1325 (mult_9_n1325, mult_9_n1376, mult_9_n13);
	xnor gate_mult_9_n1324 (mult_9_n1324, mult_9_n1375, mult_9_n13);
	xnor gate_mult_9_n1323 (mult_9_n1323, mult_9_n1374, mult_9_n13);
	xnor gate_mult_9_n1322 (mult_9_n1322, mult_9_n1373, mult_9_n13);
	xnor gate_mult_9_n1321 (mult_9_n1321, mult_9_n1372, mult_9_n13);
	xnor gate_mult_9_n1320 (mult_9_n1320, mult_9_n1371, mult_9_n13);
	xnor gate_mult_9_n1319 (mult_9_n1319, mult_9_n1370, mult_9_n13);
	xnor gate_mult_9_n1318 (mult_9_n1318, mult_9_n1369, mult_9_n13);
	xnor gate_mult_9_n1317 (mult_9_n1317, mult_9_n1368, mult_9_n13);
	xnor gate_mult_9_n1316 (mult_9_n1316, mult_9_n1367, mult_9_n13);
	xnor gate_mult_9_n1315 (mult_9_n1315, mult_9_n1366, mult_9_n13);
	xnor gate_mult_9_n1314 (mult_9_n1314, mult_9_n1365, mult_9_n13);
	xnor gate_mult_9_n1313 (mult_9_n1313, mult_9_n1364, mult_9_n13);
	xnor gate_mult_9_n1312 (mult_9_n1312, mult_9_n1363, mult_9_n13);
	not gate_mult_9_n976 (mult_9_n976, mult_9_n15);
	and gate_mult_9_n1176 (mult_9_n1176, mult_9_n49, mult_9_n976);
	or gate_mult_9_n975 (mult_9_n975, mult_9_n17, mult_9_n1327);
	or gate_mult_9_n974 (mult_9_n974, mult_9_n15, mult_9_n1326);
	nand gate_mult_9_n1175 (mult_9_n1175, mult_9_n975, mult_9_n974);
	or gate_mult_9_n973 (mult_9_n973, mult_9_n17, mult_9_n1326);
	or gate_mult_9_n972 (mult_9_n972, mult_9_n15, mult_9_n1325);
	nand gate_mult_9_n1174 (mult_9_n1174, mult_9_n973, mult_9_n972);
	or gate_mult_9_n971 (mult_9_n971, mult_9_n17, mult_9_n1325);
	or gate_mult_9_n970 (mult_9_n970, mult_9_n15, mult_9_n1324);
	nand gate_mult_9_n1173 (mult_9_n1173, mult_9_n971, mult_9_n970);
	or gate_mult_9_n969 (mult_9_n969, mult_9_n17, mult_9_n1324);
	or gate_mult_9_n968 (mult_9_n968, mult_9_n15, mult_9_n1323);
	nand gate_mult_9_n1172 (mult_9_n1172, mult_9_n969, mult_9_n968);
	or gate_mult_9_n967 (mult_9_n967, mult_9_n17, mult_9_n1323);
	or gate_mult_9_n966 (mult_9_n966, mult_9_n15, mult_9_n1322);
	nand gate_mult_9_n1171 (mult_9_n1171, mult_9_n967, mult_9_n966);
	or gate_mult_9_n965 (mult_9_n965, mult_9_n17, mult_9_n1322);
	or gate_mult_9_n964 (mult_9_n964, mult_9_n15, mult_9_n1321);
	nand gate_mult_9_n1170 (mult_9_n1170, mult_9_n965, mult_9_n964);
	or gate_mult_9_n963 (mult_9_n963, mult_9_n17, mult_9_n1321);
	or gate_mult_9_n962 (mult_9_n962, mult_9_n15, mult_9_n1320);
	nand gate_mult_9_n1169 (mult_9_n1169, mult_9_n963, mult_9_n962);
	or gate_mult_9_n961 (mult_9_n961, mult_9_n17, mult_9_n1320);
	or gate_mult_9_n960 (mult_9_n960, mult_9_n15, mult_9_n1319);
	nand gate_mult_9_n1168 (mult_9_n1168, mult_9_n961, mult_9_n960);
	or gate_mult_9_n959 (mult_9_n959, mult_9_n17, mult_9_n1319);
	or gate_mult_9_n958 (mult_9_n958, mult_9_n16, mult_9_n1318);
	nand gate_mult_9_n1167 (mult_9_n1167, mult_9_n959, mult_9_n958);
	or gate_mult_9_n957 (mult_9_n957, mult_9_n18, mult_9_n1318);
	or gate_mult_9_n956 (mult_9_n956, mult_9_n16, mult_9_n1317);
	nand gate_mult_9_n1166 (mult_9_n1166, mult_9_n957, mult_9_n956);
	or gate_mult_9_n955 (mult_9_n955, mult_9_n18, mult_9_n1317);
	or gate_mult_9_n954 (mult_9_n954, mult_9_n16, mult_9_n1316);
	nand gate_mult_9_n1165 (mult_9_n1165, mult_9_n955, mult_9_n954);
	or gate_mult_9_n953 (mult_9_n953, mult_9_n18, mult_9_n1316);
	or gate_mult_9_n952 (mult_9_n952, mult_9_n16, mult_9_n1315);
	nand gate_mult_9_n1164 (mult_9_n1164, mult_9_n953, mult_9_n952);
	or gate_mult_9_n951 (mult_9_n951, mult_9_n18, mult_9_n1315);
	or gate_mult_9_n950 (mult_9_n950, mult_9_n16, mult_9_n1314);
	nand gate_mult_9_n1163 (mult_9_n1163, mult_9_n951, mult_9_n950);
	or gate_mult_9_n949 (mult_9_n949, mult_9_n18, mult_9_n1314);
	or gate_mult_9_n948 (mult_9_n948, mult_9_n16, mult_9_n1313);
	nand gate_mult_9_n1162 (mult_9_n1162, mult_9_n949, mult_9_n948);
	or gate_mult_9_n947 (mult_9_n947, mult_9_n18, mult_9_n1313);
	or gate_mult_9_n946 (mult_9_n946, mult_9_n16, mult_9_n1312);
	nand gate_mult_9_n1161 (mult_9_n1161, mult_9_n947, mult_9_n946);
	or gate_mult_9_n945 (mult_9_n945, mult_9_n18, mult_9_n1312);
	or gate_mult_9_n944 (mult_9_n944, mult_9_n16, mult_9_n1409);
	nand gate_mult_9_n1160 (mult_9_n1160, mult_9_n945, mult_9_n944);
	and gate_mult_9_n943 (mult_9_n943, mult_9_n18, mult_9_n16);
	or gate_mult_9_n1159 (mult_9_n1159, mult_9_n1409, mult_9_n943);
	or gate_mult_9_n942 (mult_9_n942, mult_9_n16, mult_9_n1328);
	or gate_mult_9_n941 (mult_9_n941, mult_9_n18, mult_9_n1409);
	nand gate_mult_9_n1057 (mult_9_n1057, mult_9_n942, mult_9_n941);
	or gate_mult_9_n1311 (mult_9_n1311, mult_9_n49, mult_9_n1408);
	xnor gate_mult_9_n1310 (mult_9_n1310, mult_9_n49, mult_9_n19);
	xnor gate_mult_9_n1309 (mult_9_n1309, mult_9_n1377, mult_9_n19);
	xnor gate_mult_9_n1308 (mult_9_n1308, mult_9_n1376, mult_9_n19);
	xnor gate_mult_9_n1307 (mult_9_n1307, mult_9_n1375, mult_9_n19);
	xnor gate_mult_9_n1306 (mult_9_n1306, mult_9_n1374, mult_9_n19);
	xnor gate_mult_9_n1305 (mult_9_n1305, mult_9_n1373, mult_9_n19);
	xnor gate_mult_9_n1304 (mult_9_n1304, mult_9_n1372, mult_9_n19);
	xnor gate_mult_9_n1303 (mult_9_n1303, mult_9_n1371, mult_9_n19);
	xnor gate_mult_9_n1302 (mult_9_n1302, mult_9_n1370, mult_9_n19);
	xnor gate_mult_9_n1301 (mult_9_n1301, mult_9_n1369, mult_9_n19);
	xnor gate_mult_9_n1300 (mult_9_n1300, mult_9_n1368, mult_9_n19);
	xnor gate_mult_9_n1299 (mult_9_n1299, mult_9_n1367, mult_9_n19);
	xnor gate_mult_9_n1298 (mult_9_n1298, mult_9_n1366, mult_9_n19);
	xnor gate_mult_9_n1297 (mult_9_n1297, mult_9_n1365, mult_9_n19);
	xnor gate_mult_9_n1296 (mult_9_n1296, mult_9_n1364, mult_9_n19);
	xnor gate_mult_9_n1295 (mult_9_n1295, mult_9_n1363, mult_9_n19);
	not gate_mult_9_n939 (mult_9_n939, mult_9_n21);
	and gate_mult_9_n1158 (mult_9_n1158, mult_9_n49, mult_9_n939);
	or gate_mult_9_n938 (mult_9_n938, mult_9_n23, mult_9_n1310);
	or gate_mult_9_n937 (mult_9_n937, mult_9_n21, mult_9_n1309);
	nand gate_mult_9_n1157 (mult_9_n1157, mult_9_n938, mult_9_n937);
	or gate_mult_9_n936 (mult_9_n936, mult_9_n23, mult_9_n1309);
	or gate_mult_9_n935 (mult_9_n935, mult_9_n21, mult_9_n1308);
	nand gate_mult_9_n1156 (mult_9_n1156, mult_9_n936, mult_9_n935);
	or gate_mult_9_n934 (mult_9_n934, mult_9_n23, mult_9_n1308);
	or gate_mult_9_n933 (mult_9_n933, mult_9_n21, mult_9_n1307);
	nand gate_mult_9_n1155 (mult_9_n1155, mult_9_n934, mult_9_n933);
	or gate_mult_9_n932 (mult_9_n932, mult_9_n23, mult_9_n1307);
	or gate_mult_9_n931 (mult_9_n931, mult_9_n21, mult_9_n1306);
	nand gate_mult_9_n1154 (mult_9_n1154, mult_9_n932, mult_9_n931);
	or gate_mult_9_n930 (mult_9_n930, mult_9_n23, mult_9_n1306);
	or gate_mult_9_n929 (mult_9_n929, mult_9_n21, mult_9_n1305);
	nand gate_mult_9_n1153 (mult_9_n1153, mult_9_n930, mult_9_n929);
	or gate_mult_9_n928 (mult_9_n928, mult_9_n23, mult_9_n1305);
	or gate_mult_9_n927 (mult_9_n927, mult_9_n21, mult_9_n1304);
	nand gate_mult_9_n1152 (mult_9_n1152, mult_9_n928, mult_9_n927);
	or gate_mult_9_n926 (mult_9_n926, mult_9_n23, mult_9_n1304);
	or gate_mult_9_n925 (mult_9_n925, mult_9_n21, mult_9_n1303);
	nand gate_mult_9_n1151 (mult_9_n1151, mult_9_n926, mult_9_n925);
	or gate_mult_9_n924 (mult_9_n924, mult_9_n23, mult_9_n1303);
	or gate_mult_9_n923 (mult_9_n923, mult_9_n21, mult_9_n1302);
	nand gate_mult_9_n1150 (mult_9_n1150, mult_9_n924, mult_9_n923);
	or gate_mult_9_n922 (mult_9_n922, mult_9_n23, mult_9_n1302);
	or gate_mult_9_n921 (mult_9_n921, mult_9_n22, mult_9_n1301);
	nand gate_mult_9_n1149 (mult_9_n1149, mult_9_n922, mult_9_n921);
	or gate_mult_9_n920 (mult_9_n920, mult_9_n24, mult_9_n1301);
	or gate_mult_9_n919 (mult_9_n919, mult_9_n22, mult_9_n1300);
	nand gate_mult_9_n1148 (mult_9_n1148, mult_9_n920, mult_9_n919);
	or gate_mult_9_n918 (mult_9_n918, mult_9_n24, mult_9_n1300);
	or gate_mult_9_n917 (mult_9_n917, mult_9_n22, mult_9_n1299);
	nand gate_mult_9_n1147 (mult_9_n1147, mult_9_n918, mult_9_n917);
	or gate_mult_9_n916 (mult_9_n916, mult_9_n24, mult_9_n1299);
	or gate_mult_9_n915 (mult_9_n915, mult_9_n22, mult_9_n1298);
	nand gate_mult_9_n1146 (mult_9_n1146, mult_9_n916, mult_9_n915);
	or gate_mult_9_n914 (mult_9_n914, mult_9_n24, mult_9_n1298);
	or gate_mult_9_n913 (mult_9_n913, mult_9_n22, mult_9_n1297);
	nand gate_mult_9_n1145 (mult_9_n1145, mult_9_n914, mult_9_n913);
	or gate_mult_9_n912 (mult_9_n912, mult_9_n24, mult_9_n1297);
	or gate_mult_9_n911 (mult_9_n911, mult_9_n22, mult_9_n1296);
	nand gate_mult_9_n1144 (mult_9_n1144, mult_9_n912, mult_9_n911);
	or gate_mult_9_n910 (mult_9_n910, mult_9_n24, mult_9_n1296);
	or gate_mult_9_n909 (mult_9_n909, mult_9_n22, mult_9_n1295);
	nand gate_mult_9_n1143 (mult_9_n1143, mult_9_n910, mult_9_n909);
	or gate_mult_9_n908 (mult_9_n908, mult_9_n24, mult_9_n1295);
	or gate_mult_9_n907 (mult_9_n907, mult_9_n22, mult_9_n1408);
	nand gate_mult_9_n1142 (mult_9_n1142, mult_9_n908, mult_9_n907);
	and gate_mult_9_n906 (mult_9_n906, mult_9_n24, mult_9_n22);
	or gate_mult_9_n1141 (mult_9_n1141, mult_9_n1408, mult_9_n906);
	or gate_mult_9_n905 (mult_9_n905, mult_9_n22, mult_9_n1311);
	or gate_mult_9_n904 (mult_9_n904, mult_9_n24, mult_9_n1408);
	nand gate_mult_9_n1056 (mult_9_n1056, mult_9_n905, mult_9_n904);
	or gate_mult_9_n1294 (mult_9_n1294, mult_9_n49, mult_9_n1407);
	xnor gate_mult_9_n1293 (mult_9_n1293, mult_9_n49, mult_9_n25);
	xnor gate_mult_9_n1292 (mult_9_n1292, mult_9_n1377, mult_9_n25);
	xnor gate_mult_9_n1291 (mult_9_n1291, mult_9_n1376, mult_9_n25);
	xnor gate_mult_9_n1290 (mult_9_n1290, mult_9_n1375, mult_9_n25);
	xnor gate_mult_9_n1289 (mult_9_n1289, mult_9_n1374, mult_9_n25);
	xnor gate_mult_9_n1288 (mult_9_n1288, mult_9_n1373, mult_9_n25);
	xnor gate_mult_9_n1287 (mult_9_n1287, mult_9_n1372, mult_9_n25);
	xnor gate_mult_9_n1286 (mult_9_n1286, mult_9_n1371, mult_9_n25);
	xnor gate_mult_9_n1285 (mult_9_n1285, mult_9_n1370, mult_9_n25);
	xnor gate_mult_9_n1284 (mult_9_n1284, mult_9_n1369, mult_9_n25);
	xnor gate_mult_9_n1283 (mult_9_n1283, mult_9_n1368, mult_9_n25);
	xnor gate_mult_9_n1282 (mult_9_n1282, mult_9_n1367, mult_9_n25);
	xnor gate_mult_9_n1281 (mult_9_n1281, mult_9_n1366, mult_9_n25);
	xnor gate_mult_9_n1280 (mult_9_n1280, mult_9_n1365, mult_9_n25);
	xnor gate_mult_9_n1279 (mult_9_n1279, mult_9_n1364, mult_9_n25);
	xnor gate_mult_9_n1278 (mult_9_n1278, mult_9_n1363, mult_9_n25);
	not gate_mult_9_n902 (mult_9_n902, mult_9_n27);
	and gate_mult_9_n1140 (mult_9_n1140, mult_9_n49, mult_9_n902);
	or gate_mult_9_n901 (mult_9_n901, mult_9_n29, mult_9_n1293);
	or gate_mult_9_n900 (mult_9_n900, mult_9_n27, mult_9_n1292);
	nand gate_mult_9_n1139 (mult_9_n1139, mult_9_n901, mult_9_n900);
	or gate_mult_9_n899 (mult_9_n899, mult_9_n29, mult_9_n1292);
	or gate_mult_9_n898 (mult_9_n898, mult_9_n27, mult_9_n1291);
	nand gate_mult_9_n1138 (mult_9_n1138, mult_9_n899, mult_9_n898);
	or gate_mult_9_n897 (mult_9_n897, mult_9_n29, mult_9_n1291);
	or gate_mult_9_n896 (mult_9_n896, mult_9_n27, mult_9_n1290);
	nand gate_mult_9_n1137 (mult_9_n1137, mult_9_n897, mult_9_n896);
	or gate_mult_9_n895 (mult_9_n895, mult_9_n29, mult_9_n1290);
	or gate_mult_9_n894 (mult_9_n894, mult_9_n27, mult_9_n1289);
	nand gate_mult_9_n1136 (mult_9_n1136, mult_9_n895, mult_9_n894);
	or gate_mult_9_n893 (mult_9_n893, mult_9_n29, mult_9_n1289);
	or gate_mult_9_n892 (mult_9_n892, mult_9_n27, mult_9_n1288);
	nand gate_mult_9_n1135 (mult_9_n1135, mult_9_n893, mult_9_n892);
	or gate_mult_9_n891 (mult_9_n891, mult_9_n29, mult_9_n1288);
	or gate_mult_9_n890 (mult_9_n890, mult_9_n27, mult_9_n1287);
	nand gate_mult_9_n1134 (mult_9_n1134, mult_9_n891, mult_9_n890);
	or gate_mult_9_n889 (mult_9_n889, mult_9_n29, mult_9_n1287);
	or gate_mult_9_n888 (mult_9_n888, mult_9_n27, mult_9_n1286);
	nand gate_mult_9_n1133 (mult_9_n1133, mult_9_n889, mult_9_n888);
	or gate_mult_9_n887 (mult_9_n887, mult_9_n29, mult_9_n1286);
	or gate_mult_9_n886 (mult_9_n886, mult_9_n27, mult_9_n1285);
	nand gate_mult_9_n1132 (mult_9_n1132, mult_9_n887, mult_9_n886);
	or gate_mult_9_n885 (mult_9_n885, mult_9_n29, mult_9_n1285);
	or gate_mult_9_n884 (mult_9_n884, mult_9_n28, mult_9_n1284);
	nand gate_mult_9_n1131 (mult_9_n1131, mult_9_n885, mult_9_n884);
	or gate_mult_9_n883 (mult_9_n883, mult_9_n30, mult_9_n1284);
	or gate_mult_9_n882 (mult_9_n882, mult_9_n28, mult_9_n1283);
	nand gate_mult_9_n1130 (mult_9_n1130, mult_9_n883, mult_9_n882);
	or gate_mult_9_n881 (mult_9_n881, mult_9_n30, mult_9_n1283);
	or gate_mult_9_n880 (mult_9_n880, mult_9_n28, mult_9_n1282);
	nand gate_mult_9_n1129 (mult_9_n1129, mult_9_n881, mult_9_n880);
	or gate_mult_9_n879 (mult_9_n879, mult_9_n30, mult_9_n1282);
	or gate_mult_9_n878 (mult_9_n878, mult_9_n28, mult_9_n1281);
	nand gate_mult_9_n1128 (mult_9_n1128, mult_9_n879, mult_9_n878);
	or gate_mult_9_n877 (mult_9_n877, mult_9_n30, mult_9_n1281);
	or gate_mult_9_n876 (mult_9_n876, mult_9_n28, mult_9_n1280);
	nand gate_mult_9_n1127 (mult_9_n1127, mult_9_n877, mult_9_n876);
	or gate_mult_9_n875 (mult_9_n875, mult_9_n30, mult_9_n1280);
	or gate_mult_9_n874 (mult_9_n874, mult_9_n28, mult_9_n1279);
	nand gate_mult_9_n1126 (mult_9_n1126, mult_9_n875, mult_9_n874);
	or gate_mult_9_n873 (mult_9_n873, mult_9_n30, mult_9_n1279);
	or gate_mult_9_n872 (mult_9_n872, mult_9_n28, mult_9_n1278);
	nand gate_mult_9_n1125 (mult_9_n1125, mult_9_n873, mult_9_n872);
	or gate_mult_9_n871 (mult_9_n871, mult_9_n30, mult_9_n1278);
	or gate_mult_9_n870 (mult_9_n870, mult_9_n28, mult_9_n1407);
	nand gate_mult_9_n1124 (mult_9_n1124, mult_9_n871, mult_9_n870);
	and gate_mult_9_n869 (mult_9_n869, mult_9_n30, mult_9_n28);
	or gate_mult_9_n1123 (mult_9_n1123, mult_9_n1407, mult_9_n869);
	or gate_mult_9_n868 (mult_9_n868, mult_9_n28, mult_9_n1294);
	or gate_mult_9_n867 (mult_9_n867, mult_9_n30, mult_9_n1407);
	nand gate_mult_9_n1055 (mult_9_n1055, mult_9_n868, mult_9_n867);
	or gate_mult_9_n1277 (mult_9_n1277, mult_9_n49, mult_9_n1406);
	xnor gate_mult_9_n1276 (mult_9_n1276, mult_9_n49, mult_9_n31);
	xnor gate_mult_9_n1275 (mult_9_n1275, mult_9_n1377, mult_9_n31);
	xnor gate_mult_9_n1274 (mult_9_n1274, mult_9_n1376, mult_9_n31);
	xnor gate_mult_9_n1273 (mult_9_n1273, mult_9_n1375, mult_9_n31);
	xnor gate_mult_9_n1272 (mult_9_n1272, mult_9_n1374, mult_9_n31);
	xnor gate_mult_9_n1271 (mult_9_n1271, mult_9_n1373, mult_9_n31);
	xnor gate_mult_9_n1270 (mult_9_n1270, mult_9_n1372, mult_9_n31);
	xnor gate_mult_9_n1269 (mult_9_n1269, mult_9_n1371, mult_9_n31);
	xnor gate_mult_9_n1268 (mult_9_n1268, mult_9_n1370, mult_9_n31);
	xnor gate_mult_9_n1267 (mult_9_n1267, mult_9_n1369, mult_9_n31);
	xnor gate_mult_9_n1266 (mult_9_n1266, mult_9_n1368, mult_9_n31);
	xnor gate_mult_9_n1265 (mult_9_n1265, mult_9_n1367, mult_9_n31);
	xnor gate_mult_9_n1264 (mult_9_n1264, mult_9_n1366, mult_9_n31);
	xnor gate_mult_9_n1263 (mult_9_n1263, mult_9_n1365, mult_9_n31);
	xnor gate_mult_9_n1262 (mult_9_n1262, mult_9_n1364, mult_9_n31);
	xnor gate_mult_9_n1261 (mult_9_n1261, mult_9_n1363, mult_9_n31);
	not gate_mult_9_n865 (mult_9_n865, mult_9_n33);
	and gate_mult_9_n1122 (mult_9_n1122, mult_9_n49, mult_9_n865);
	or gate_mult_9_n864 (mult_9_n864, mult_9_n35, mult_9_n1276);
	or gate_mult_9_n863 (mult_9_n863, mult_9_n33, mult_9_n1275);
	nand gate_mult_9_n1121 (mult_9_n1121, mult_9_n864, mult_9_n863);
	or gate_mult_9_n862 (mult_9_n862, mult_9_n35, mult_9_n1275);
	or gate_mult_9_n861 (mult_9_n861, mult_9_n33, mult_9_n1274);
	nand gate_mult_9_n1120 (mult_9_n1120, mult_9_n862, mult_9_n861);
	or gate_mult_9_n860 (mult_9_n860, mult_9_n35, mult_9_n1274);
	or gate_mult_9_n859 (mult_9_n859, mult_9_n33, mult_9_n1273);
	nand gate_mult_9_n1119 (mult_9_n1119, mult_9_n860, mult_9_n859);
	or gate_mult_9_n858 (mult_9_n858, mult_9_n35, mult_9_n1273);
	or gate_mult_9_n857 (mult_9_n857, mult_9_n33, mult_9_n1272);
	nand gate_mult_9_n1118 (mult_9_n1118, mult_9_n858, mult_9_n857);
	or gate_mult_9_n856 (mult_9_n856, mult_9_n35, mult_9_n1272);
	or gate_mult_9_n855 (mult_9_n855, mult_9_n33, mult_9_n1271);
	nand gate_mult_9_n1117 (mult_9_n1117, mult_9_n856, mult_9_n855);
	or gate_mult_9_n854 (mult_9_n854, mult_9_n35, mult_9_n1271);
	or gate_mult_9_n853 (mult_9_n853, mult_9_n33, mult_9_n1270);
	nand gate_mult_9_n1116 (mult_9_n1116, mult_9_n854, mult_9_n853);
	or gate_mult_9_n852 (mult_9_n852, mult_9_n35, mult_9_n1270);
	or gate_mult_9_n851 (mult_9_n851, mult_9_n33, mult_9_n1269);
	nand gate_mult_9_n1115 (mult_9_n1115, mult_9_n852, mult_9_n851);
	or gate_mult_9_n850 (mult_9_n850, mult_9_n35, mult_9_n1269);
	or gate_mult_9_n849 (mult_9_n849, mult_9_n33, mult_9_n1268);
	nand gate_mult_9_n1114 (mult_9_n1114, mult_9_n850, mult_9_n849);
	or gate_mult_9_n848 (mult_9_n848, mult_9_n35, mult_9_n1268);
	or gate_mult_9_n847 (mult_9_n847, mult_9_n34, mult_9_n1267);
	nand gate_mult_9_n1113 (mult_9_n1113, mult_9_n848, mult_9_n847);
	or gate_mult_9_n846 (mult_9_n846, mult_9_n36, mult_9_n1267);
	or gate_mult_9_n845 (mult_9_n845, mult_9_n34, mult_9_n1266);
	nand gate_mult_9_n1112 (mult_9_n1112, mult_9_n846, mult_9_n845);
	or gate_mult_9_n844 (mult_9_n844, mult_9_n36, mult_9_n1266);
	or gate_mult_9_n843 (mult_9_n843, mult_9_n34, mult_9_n1265);
	nand gate_mult_9_n1111 (mult_9_n1111, mult_9_n844, mult_9_n843);
	or gate_mult_9_n842 (mult_9_n842, mult_9_n36, mult_9_n1265);
	or gate_mult_9_n841 (mult_9_n841, mult_9_n34, mult_9_n1264);
	nand gate_mult_9_n1110 (mult_9_n1110, mult_9_n842, mult_9_n841);
	or gate_mult_9_n840 (mult_9_n840, mult_9_n36, mult_9_n1264);
	or gate_mult_9_n839 (mult_9_n839, mult_9_n34, mult_9_n1263);
	nand gate_mult_9_n1109 (mult_9_n1109, mult_9_n840, mult_9_n839);
	or gate_mult_9_n838 (mult_9_n838, mult_9_n36, mult_9_n1263);
	or gate_mult_9_n837 (mult_9_n837, mult_9_n34, mult_9_n1262);
	nand gate_mult_9_n1108 (mult_9_n1108, mult_9_n838, mult_9_n837);
	or gate_mult_9_n836 (mult_9_n836, mult_9_n36, mult_9_n1262);
	or gate_mult_9_n835 (mult_9_n835, mult_9_n34, mult_9_n1261);
	nand gate_mult_9_n1107 (mult_9_n1107, mult_9_n836, mult_9_n835);
	or gate_mult_9_n834 (mult_9_n834, mult_9_n36, mult_9_n1261);
	or gate_mult_9_n833 (mult_9_n833, mult_9_n34, mult_9_n1406);
	nand gate_mult_9_n1106 (mult_9_n1106, mult_9_n834, mult_9_n833);
	and gate_mult_9_n832 (mult_9_n832, mult_9_n36, mult_9_n34);
	or gate_mult_9_n1105 (mult_9_n1105, mult_9_n1406, mult_9_n832);
	or gate_mult_9_n831 (mult_9_n831, mult_9_n34, mult_9_n1277);
	or gate_mult_9_n830 (mult_9_n830, mult_9_n36, mult_9_n1406);
	nand gate_mult_9_n1054 (mult_9_n1054, mult_9_n831, mult_9_n830);
	or gate_mult_9_n1260 (mult_9_n1260, mult_9_n49, mult_9_n1405);
	xnor gate_mult_9_n1259 (mult_9_n1259, mult_9_n49, mult_9_n37);
	xnor gate_mult_9_n1258 (mult_9_n1258, mult_9_n1377, mult_9_n37);
	xnor gate_mult_9_n1257 (mult_9_n1257, mult_9_n1376, mult_9_n37);
	xnor gate_mult_9_n1256 (mult_9_n1256, mult_9_n1375, mult_9_n37);
	xnor gate_mult_9_n1255 (mult_9_n1255, mult_9_n1374, mult_9_n37);
	xnor gate_mult_9_n1254 (mult_9_n1254, mult_9_n1373, mult_9_n37);
	xnor gate_mult_9_n1253 (mult_9_n1253, mult_9_n1372, mult_9_n37);
	xnor gate_mult_9_n1252 (mult_9_n1252, mult_9_n1371, mult_9_n37);
	xnor gate_mult_9_n1251 (mult_9_n1251, mult_9_n1370, mult_9_n37);
	xnor gate_mult_9_n1250 (mult_9_n1250, mult_9_n1369, mult_9_n37);
	xnor gate_mult_9_n1249 (mult_9_n1249, mult_9_n1368, mult_9_n37);
	xnor gate_mult_9_n1248 (mult_9_n1248, mult_9_n1367, mult_9_n37);
	xnor gate_mult_9_n1247 (mult_9_n1247, mult_9_n1366, mult_9_n37);
	xnor gate_mult_9_n1246 (mult_9_n1246, mult_9_n1365, mult_9_n37);
	xnor gate_mult_9_n1245 (mult_9_n1245, mult_9_n1364, mult_9_n37);
	xnor gate_mult_9_n1244 (mult_9_n1244, mult_9_n1363, mult_9_n37);
	not gate_mult_9_n828 (mult_9_n828, mult_9_n39);
	and gate_mult_9_n1104 (mult_9_n1104, mult_9_n49, mult_9_n828);
	or gate_mult_9_n827 (mult_9_n827, mult_9_n41, mult_9_n1259);
	or gate_mult_9_n826 (mult_9_n826, mult_9_n39, mult_9_n1258);
	nand gate_mult_9_n1103 (mult_9_n1103, mult_9_n827, mult_9_n826);
	or gate_mult_9_n825 (mult_9_n825, mult_9_n41, mult_9_n1258);
	or gate_mult_9_n824 (mult_9_n824, mult_9_n39, mult_9_n1257);
	nand gate_mult_9_n1102 (mult_9_n1102, mult_9_n825, mult_9_n824);
	or gate_mult_9_n823 (mult_9_n823, mult_9_n41, mult_9_n1257);
	or gate_mult_9_n822 (mult_9_n822, mult_9_n39, mult_9_n1256);
	nand gate_mult_9_n1101 (mult_9_n1101, mult_9_n823, mult_9_n822);
	or gate_mult_9_n821 (mult_9_n821, mult_9_n41, mult_9_n1256);
	or gate_mult_9_n820 (mult_9_n820, mult_9_n39, mult_9_n1255);
	nand gate_mult_9_n1100 (mult_9_n1100, mult_9_n821, mult_9_n820);
	or gate_mult_9_n819 (mult_9_n819, mult_9_n41, mult_9_n1255);
	or gate_mult_9_n818 (mult_9_n818, mult_9_n39, mult_9_n1254);
	nand gate_mult_9_n1099 (mult_9_n1099, mult_9_n819, mult_9_n818);
	or gate_mult_9_n817 (mult_9_n817, mult_9_n41, mult_9_n1254);
	or gate_mult_9_n816 (mult_9_n816, mult_9_n39, mult_9_n1253);
	nand gate_mult_9_n1098 (mult_9_n1098, mult_9_n817, mult_9_n816);
	or gate_mult_9_n815 (mult_9_n815, mult_9_n41, mult_9_n1253);
	or gate_mult_9_n814 (mult_9_n814, mult_9_n39, mult_9_n1252);
	nand gate_mult_9_n1097 (mult_9_n1097, mult_9_n815, mult_9_n814);
	or gate_mult_9_n813 (mult_9_n813, mult_9_n41, mult_9_n1252);
	or gate_mult_9_n812 (mult_9_n812, mult_9_n39, mult_9_n1251);
	nand gate_mult_9_n1096 (mult_9_n1096, mult_9_n813, mult_9_n812);
	or gate_mult_9_n811 (mult_9_n811, mult_9_n41, mult_9_n1251);
	or gate_mult_9_n810 (mult_9_n810, mult_9_n40, mult_9_n1250);
	nand gate_mult_9_n1095 (mult_9_n1095, mult_9_n811, mult_9_n810);
	or gate_mult_9_n809 (mult_9_n809, mult_9_n42, mult_9_n1250);
	or gate_mult_9_n808 (mult_9_n808, mult_9_n40, mult_9_n1249);
	nand gate_mult_9_n1094 (mult_9_n1094, mult_9_n809, mult_9_n808);
	or gate_mult_9_n807 (mult_9_n807, mult_9_n42, mult_9_n1249);
	or gate_mult_9_n806 (mult_9_n806, mult_9_n40, mult_9_n1248);
	nand gate_mult_9_n1093 (mult_9_n1093, mult_9_n807, mult_9_n806);
	or gate_mult_9_n805 (mult_9_n805, mult_9_n42, mult_9_n1248);
	or gate_mult_9_n804 (mult_9_n804, mult_9_n40, mult_9_n1247);
	nand gate_mult_9_n1092 (mult_9_n1092, mult_9_n805, mult_9_n804);
	or gate_mult_9_n803 (mult_9_n803, mult_9_n42, mult_9_n1247);
	or gate_mult_9_n802 (mult_9_n802, mult_9_n40, mult_9_n1246);
	nand gate_mult_9_n1091 (mult_9_n1091, mult_9_n803, mult_9_n802);
	or gate_mult_9_n801 (mult_9_n801, mult_9_n42, mult_9_n1246);
	or gate_mult_9_n800 (mult_9_n800, mult_9_n40, mult_9_n1245);
	nand gate_mult_9_n1090 (mult_9_n1090, mult_9_n801, mult_9_n800);
	or gate_mult_9_n799 (mult_9_n799, mult_9_n42, mult_9_n1245);
	or gate_mult_9_n798 (mult_9_n798, mult_9_n40, mult_9_n1244);
	nand gate_mult_9_n1089 (mult_9_n1089, mult_9_n799, mult_9_n798);
	or gate_mult_9_n797 (mult_9_n797, mult_9_n42, mult_9_n1244);
	or gate_mult_9_n796 (mult_9_n796, mult_9_n40, mult_9_n1405);
	nand gate_mult_9_n1088 (mult_9_n1088, mult_9_n797, mult_9_n796);
	and gate_mult_9_n795 (mult_9_n795, mult_9_n42, mult_9_n40);
	or gate_mult_9_n1087 (mult_9_n1087, mult_9_n1405, mult_9_n795);
	or gate_mult_9_n794 (mult_9_n794, mult_9_n40, mult_9_n1260);
	or gate_mult_9_n793 (mult_9_n793, mult_9_n42, mult_9_n1405);
	nand gate_mult_9_n1053 (mult_9_n1053, mult_9_n794, mult_9_n793);
	or gate_mult_9_n1243 (mult_9_n1243, mult_9_n49, mult_9_n1404);
	xnor gate_mult_9_n1242 (mult_9_n1242, mult_9_n49, mult_9_n43);
	xnor gate_mult_9_n1241 (mult_9_n1241, mult_9_n1377, mult_9_n43);
	xnor gate_mult_9_n1240 (mult_9_n1240, mult_9_n1376, mult_9_n43);
	xnor gate_mult_9_n1239 (mult_9_n1239, mult_9_n1375, mult_9_n43);
	xnor gate_mult_9_n1238 (mult_9_n1238, mult_9_n1374, mult_9_n43);
	xnor gate_mult_9_n1237 (mult_9_n1237, mult_9_n1373, mult_9_n43);
	xnor gate_mult_9_n1236 (mult_9_n1236, mult_9_n1372, mult_9_n43);
	xnor gate_mult_9_n1235 (mult_9_n1235, mult_9_n1371, mult_9_n43);
	xnor gate_mult_9_n1234 (mult_9_n1234, mult_9_n1370, mult_9_n43);
	xnor gate_mult_9_n1233 (mult_9_n1233, mult_9_n1369, mult_9_n43);
	xnor gate_mult_9_n1232 (mult_9_n1232, mult_9_n1368, mult_9_n43);
	xnor gate_mult_9_n1231 (mult_9_n1231, mult_9_n1367, mult_9_n43);
	xnor gate_mult_9_n1230 (mult_9_n1230, mult_9_n1366, mult_9_n43);
	xnor gate_mult_9_n1229 (mult_9_n1229, mult_9_n1365, mult_9_n43);
	xnor gate_mult_9_n1228 (mult_9_n1228, mult_9_n1364, mult_9_n43);
	xnor gate_mult_9_n1227 (mult_9_n1227, mult_9_n1363, mult_9_n43);
	not gate_mult_9_n791 (mult_9_n791, mult_9_n45);
	and gate_mult_9_n1086 (mult_9_n1086, mult_9_n49, mult_9_n791);
	or gate_mult_9_n790 (mult_9_n790, mult_9_n47, mult_9_n1242);
	or gate_mult_9_n789 (mult_9_n789, mult_9_n45, mult_9_n1241);
	nand gate_mult_9_n1085 (mult_9_n1085, mult_9_n790, mult_9_n789);
	or gate_mult_9_n788 (mult_9_n788, mult_9_n47, mult_9_n1241);
	or gate_mult_9_n787 (mult_9_n787, mult_9_n45, mult_9_n1240);
	nand gate_mult_9_n1084 (mult_9_n1084, mult_9_n788, mult_9_n787);
	or gate_mult_9_n786 (mult_9_n786, mult_9_n47, mult_9_n1240);
	or gate_mult_9_n785 (mult_9_n785, mult_9_n45, mult_9_n1239);
	nand gate_mult_9_n1083 (mult_9_n1083, mult_9_n786, mult_9_n785);
	or gate_mult_9_n784 (mult_9_n784, mult_9_n47, mult_9_n1239);
	or gate_mult_9_n783 (mult_9_n783, mult_9_n45, mult_9_n1238);
	nand gate_mult_9_n1082 (mult_9_n1082, mult_9_n784, mult_9_n783);
	or gate_mult_9_n782 (mult_9_n782, mult_9_n47, mult_9_n1238);
	or gate_mult_9_n781 (mult_9_n781, mult_9_n45, mult_9_n1237);
	nand gate_mult_9_n1081 (mult_9_n1081, mult_9_n782, mult_9_n781);
	or gate_mult_9_n780 (mult_9_n780, mult_9_n47, mult_9_n1237);
	or gate_mult_9_n779 (mult_9_n779, mult_9_n45, mult_9_n1236);
	nand gate_mult_9_n1080 (mult_9_n1080, mult_9_n780, mult_9_n779);
	or gate_mult_9_n778 (mult_9_n778, mult_9_n47, mult_9_n1236);
	or gate_mult_9_n777 (mult_9_n777, mult_9_n45, mult_9_n1235);
	nand gate_mult_9_n1079 (mult_9_n1079, mult_9_n778, mult_9_n777);
	or gate_mult_9_n776 (mult_9_n776, mult_9_n47, mult_9_n1235);
	or gate_mult_9_n775 (mult_9_n775, mult_9_n45, mult_9_n1234);
	nand gate_mult_9_n1078 (mult_9_n1078, mult_9_n776, mult_9_n775);
	or gate_mult_9_n774 (mult_9_n774, mult_9_n47, mult_9_n1234);
	or gate_mult_9_n773 (mult_9_n773, mult_9_n46, mult_9_n1233);
	nand gate_mult_9_n1077 (mult_9_n1077, mult_9_n774, mult_9_n773);
	or gate_mult_9_n772 (mult_9_n772, mult_9_n48, mult_9_n1233);
	or gate_mult_9_n771 (mult_9_n771, mult_9_n46, mult_9_n1232);
	nand gate_mult_9_n1076 (mult_9_n1076, mult_9_n772, mult_9_n771);
	or gate_mult_9_n770 (mult_9_n770, mult_9_n48, mult_9_n1232);
	or gate_mult_9_n769 (mult_9_n769, mult_9_n46, mult_9_n1231);
	nand gate_mult_9_n1075 (mult_9_n1075, mult_9_n770, mult_9_n769);
	or gate_mult_9_n768 (mult_9_n768, mult_9_n48, mult_9_n1231);
	or gate_mult_9_n767 (mult_9_n767, mult_9_n46, mult_9_n1230);
	nand gate_mult_9_n1074 (mult_9_n1074, mult_9_n768, mult_9_n767);
	or gate_mult_9_n766 (mult_9_n766, mult_9_n48, mult_9_n1230);
	or gate_mult_9_n765 (mult_9_n765, mult_9_n46, mult_9_n1229);
	nand gate_mult_9_n1073 (mult_9_n1073, mult_9_n766, mult_9_n765);
	or gate_mult_9_n764 (mult_9_n764, mult_9_n48, mult_9_n1229);
	or gate_mult_9_n763 (mult_9_n763, mult_9_n46, mult_9_n1228);
	nand gate_mult_9_n1072 (mult_9_n1072, mult_9_n764, mult_9_n763);
	or gate_mult_9_n762 (mult_9_n762, mult_9_n48, mult_9_n1228);
	or gate_mult_9_n761 (mult_9_n761, mult_9_n46, mult_9_n1227);
	nand gate_mult_9_n1071 (mult_9_n1071, mult_9_n762, mult_9_n761);
	or gate_mult_9_n760 (mult_9_n760, mult_9_n48, mult_9_n1227);
	or gate_mult_9_n759 (mult_9_n759, mult_9_n46, mult_9_n1404);
	nand gate_mult_9_n1070 (mult_9_n1070, mult_9_n760, mult_9_n759);
	and gate_mult_9_n758 (mult_9_n758, mult_9_n48, mult_9_n46);
	or gate_mult_9_n1069 (mult_9_n1069, mult_9_n1404, mult_9_n758);
	or gate_mult_9_n757 (mult_9_n757, mult_9_n46, mult_9_n1243);
	or gate_mult_9_n756 (mult_9_n756, mult_9_n48, mult_9_n1404);
	nand gate_mult_9_n1052 (mult_9_n1052, mult_9_n757, mult_9_n756);
	not gate_mult_9_n1226 (mult_9_n1226, mult_9_n1377);
	not gate_mult_9_n1225 (mult_9_n1225, mult_9_n1376);
	not gate_mult_9_n1224 (mult_9_n1224, mult_9_n1375);
	not gate_mult_9_n1223 (mult_9_n1223, mult_9_n1374);
	not gate_mult_9_n1222 (mult_9_n1222, mult_9_n1373);
	not gate_mult_9_n1221 (mult_9_n1221, mult_9_n1372);
	not gate_mult_9_n1220 (mult_9_n1220, mult_9_n1371);
	not gate_mult_9_n1219 (mult_9_n1219, mult_9_n1370);
	not gate_mult_9_n1218 (mult_9_n1218, mult_9_n1369);
	not gate_mult_9_n1217 (mult_9_n1217, mult_9_n1368);
	not gate_mult_9_n1216 (mult_9_n1216, mult_9_n1367);
	not gate_mult_9_n1215 (mult_9_n1215, mult_9_n1366);
	not gate_mult_9_n1214 (mult_9_n1214, mult_9_n1365);
	not gate_mult_9_n1213 (mult_9_n1213, mult_9_n1364);
	not gate_mult_9_n1212 (mult_9_n1212, mult_9_n1363);
	not gate_mult_9_n755 (mult_9_n755, mult_9_n1395);
	and gate_mult_9_n1068 (mult_9_n1068, mult_9_n49, mult_9_n755);
	nor gate_mult_9_n458 (mult_9_n458, mult_9_n1226, mult_9_n1395);
	nor gate_mult_9_n1067 (mult_9_n1067, mult_9_n1225, mult_9_n1395);
	nor gate_mult_9_n1066 (mult_9_n1066, mult_9_n1224, mult_9_n1395);
	nor gate_mult_9_n386 (mult_9_n386, mult_9_n1223, mult_9_n1395);
	nor gate_mult_9_n1065 (mult_9_n1065, mult_9_n1222, mult_9_n1395);
	nor gate_mult_9_n324 (mult_9_n324, mult_9_n1221, mult_9_n1395);
	nor gate_mult_9_n1064 (mult_9_n1064, mult_9_n1220, mult_9_n1395);
	nor gate_mult_9_n272 (mult_9_n272, mult_9_n1219, mult_9_n1395);
	nor gate_mult_9_n1063 (mult_9_n1063, mult_9_n1218, mult_9_n1395);
	nor gate_mult_9_n230 (mult_9_n230, mult_9_n1217, mult_9_n1395);
	nor gate_mult_9_n1062 (mult_9_n1062, mult_9_n1216, mult_9_n1395);
	nor gate_mult_9_n198 (mult_9_n198, mult_9_n1215, mult_9_n1395);
	nor gate_mult_9_n1061 (mult_9_n1061, mult_9_n1214, mult_9_n1395);
	nor gate_mult_9_n176 (mult_9_n176, mult_9_n1213, mult_9_n1395);
	nor gate_mult_9_n1060 (mult_9_n1060, mult_9_n1212, mult_9_n1395);
	and gate_mult_9_n753 (mult_9_n753, mult_9_n1193, mult_9_n1209);
	xor gate_mult_9_n754 (mult_9_n754, mult_9_n1209, mult_9_n1193);
	xor gate_mult_9_n750 (mult_9_n750, mult_9_n1208, mult_9_n1192);
	and gate_mult_9_n749 (mult_9_n749, mult_9_n1192, mult_9_n1208);
	and gate_mult_9_n748 (mult_9_n748, mult_9_n750, mult_9_n1176);
	or gate_mult_9_n751 (mult_9_n751, mult_9_n749, mult_9_n748);
	xor gate_mult_9_n752 (mult_9_n752, mult_9_n1176, mult_9_n750);
	and gate_mult_9_n746 (mult_9_n746, mult_9_n1057, mult_9_n1207);
	xor gate_mult_9_n747 (mult_9_n747, mult_9_n1207, mult_9_n1057);
	xor gate_mult_9_n743 (mult_9_n743, mult_9_n1191, mult_9_n1175);
	and gate_mult_9_n742 (mult_9_n742, mult_9_n1175, mult_9_n1191);
	and gate_mult_9_n741 (mult_9_n741, mult_9_n747, mult_9_n743);
	or gate_mult_9_n744 (mult_9_n744, mult_9_n742, mult_9_n741);
	xor gate_mult_9_n745 (mult_9_n745, mult_9_n743, mult_9_n747);
	xor gate_mult_9_n738 (mult_9_n738, mult_9_n1206, mult_9_n1190);
	and gate_mult_9_n737 (mult_9_n737, mult_9_n1190, mult_9_n1206);
	and gate_mult_9_n736 (mult_9_n736, mult_9_n738, mult_9_n1174);
	or gate_mult_9_n739 (mult_9_n739, mult_9_n737, mult_9_n736);
	xor gate_mult_9_n740 (mult_9_n740, mult_9_n1174, mult_9_n738);
	xor gate_mult_9_n733 (mult_9_n733, mult_9_n1158, mult_9_n746);
	and gate_mult_9_n732 (mult_9_n732, mult_9_n746, mult_9_n1158);
	and gate_mult_9_n731 (mult_9_n731, mult_9_n744, mult_9_n733);
	or gate_mult_9_n734 (mult_9_n734, mult_9_n732, mult_9_n731);
	xor gate_mult_9_n735 (mult_9_n735, mult_9_n733, mult_9_n744);
	and gate_mult_9_n729 (mult_9_n729, mult_9_n1056, mult_9_n1205);
	xor gate_mult_9_n730 (mult_9_n730, mult_9_n1205, mult_9_n1056);
	xor gate_mult_9_n726 (mult_9_n726, mult_9_n1189, mult_9_n1173);
	and gate_mult_9_n725 (mult_9_n725, mult_9_n1173, mult_9_n1189);
	and gate_mult_9_n724 (mult_9_n724, mult_9_n726, mult_9_n1157);
	or gate_mult_9_n727 (mult_9_n727, mult_9_n725, mult_9_n724);
	xor gate_mult_9_n728 (mult_9_n728, mult_9_n1157, mult_9_n726);
	xor gate_mult_9_n721 (mult_9_n721, mult_9_n730, mult_9_n739);
	and gate_mult_9_n720 (mult_9_n720, mult_9_n739, mult_9_n730);
	and gate_mult_9_n719 (mult_9_n719, mult_9_n721, mult_9_n728);
	or gate_mult_9_n722 (mult_9_n722, mult_9_n720, mult_9_n719);
	xor gate_mult_9_n723 (mult_9_n723, mult_9_n728, mult_9_n721);
	xor gate_mult_9_n716 (mult_9_n716, mult_9_n1204, mult_9_n1188);
	and gate_mult_9_n715 (mult_9_n715, mult_9_n1188, mult_9_n1204);
	and gate_mult_9_n714 (mult_9_n714, mult_9_n716, mult_9_n1172);
	or gate_mult_9_n717 (mult_9_n717, mult_9_n715, mult_9_n714);
	xor gate_mult_9_n718 (mult_9_n718, mult_9_n1172, mult_9_n716);
	xor gate_mult_9_n711 (mult_9_n711, mult_9_n1156, mult_9_n1140);
	and gate_mult_9_n710 (mult_9_n710, mult_9_n1140, mult_9_n1156);
	and gate_mult_9_n709 (mult_9_n709, mult_9_n711, mult_9_n729);
	or gate_mult_9_n712 (mult_9_n712, mult_9_n710, mult_9_n709);
	xor gate_mult_9_n713 (mult_9_n713, mult_9_n729, mult_9_n711);
	xor gate_mult_9_n706 (mult_9_n706, mult_9_n727, mult_9_n718);
	and gate_mult_9_n705 (mult_9_n705, mult_9_n718, mult_9_n727);
	and gate_mult_9_n704 (mult_9_n704, mult_9_n706, mult_9_n713);
	or gate_mult_9_n707 (mult_9_n707, mult_9_n705, mult_9_n704);
	xor gate_mult_9_n708 (mult_9_n708, mult_9_n713, mult_9_n706);
	and gate_mult_9_n702 (mult_9_n702, mult_9_n1055, mult_9_n1203);
	xor gate_mult_9_n703 (mult_9_n703, mult_9_n1203, mult_9_n1055);
	xor gate_mult_9_n699 (mult_9_n699, mult_9_n1155, mult_9_n1187);
	and gate_mult_9_n698 (mult_9_n698, mult_9_n1187, mult_9_n1155);
	and gate_mult_9_n697 (mult_9_n697, mult_9_n699, mult_9_n1171);
	or gate_mult_9_n700 (mult_9_n700, mult_9_n698, mult_9_n697);
	xor gate_mult_9_n701 (mult_9_n701, mult_9_n1171, mult_9_n699);
	xor gate_mult_9_n694 (mult_9_n694, mult_9_n1139, mult_9_n703);
	and gate_mult_9_n693 (mult_9_n693, mult_9_n703, mult_9_n1139);
	and gate_mult_9_n692 (mult_9_n692, mult_9_n694, mult_9_n717);
	or gate_mult_9_n695 (mult_9_n695, mult_9_n693, mult_9_n692);
	xor gate_mult_9_n696 (mult_9_n696, mult_9_n717, mult_9_n694);
	xor gate_mult_9_n689 (mult_9_n689, mult_9_n712, mult_9_n701);
	and gate_mult_9_n688 (mult_9_n688, mult_9_n701, mult_9_n712);
	and gate_mult_9_n687 (mult_9_n687, mult_9_n696, mult_9_n689);
	or gate_mult_9_n690 (mult_9_n690, mult_9_n688, mult_9_n687);
	xor gate_mult_9_n691 (mult_9_n691, mult_9_n689, mult_9_n696);
	xor gate_mult_9_n684 (mult_9_n684, mult_9_n1202, mult_9_n1186);
	and gate_mult_9_n683 (mult_9_n683, mult_9_n1186, mult_9_n1202);
	and gate_mult_9_n682 (mult_9_n682, mult_9_n684, mult_9_n1170);
	or gate_mult_9_n685 (mult_9_n685, mult_9_n683, mult_9_n682);
	xor gate_mult_9_n686 (mult_9_n686, mult_9_n1170, mult_9_n684);
	xor gate_mult_9_n679 (mult_9_n679, mult_9_n1154, mult_9_n1138);
	and gate_mult_9_n678 (mult_9_n678, mult_9_n1138, mult_9_n1154);
	and gate_mult_9_n677 (mult_9_n677, mult_9_n679, mult_9_n1122);
	or gate_mult_9_n680 (mult_9_n680, mult_9_n678, mult_9_n677);
	xor gate_mult_9_n681 (mult_9_n681, mult_9_n1122, mult_9_n679);
	xor gate_mult_9_n674 (mult_9_n674, mult_9_n702, mult_9_n700);
	and gate_mult_9_n673 (mult_9_n673, mult_9_n700, mult_9_n702);
	and gate_mult_9_n672 (mult_9_n672, mult_9_n674, mult_9_n686);
	or gate_mult_9_n675 (mult_9_n675, mult_9_n673, mult_9_n672);
	xor gate_mult_9_n676 (mult_9_n676, mult_9_n686, mult_9_n674);
	xor gate_mult_9_n669 (mult_9_n669, mult_9_n681, mult_9_n695);
	and gate_mult_9_n668 (mult_9_n668, mult_9_n695, mult_9_n681);
	and gate_mult_9_n667 (mult_9_n667, mult_9_n676, mult_9_n669);
	or gate_mult_9_n670 (mult_9_n670, mult_9_n668, mult_9_n667);
	xor gate_mult_9_n671 (mult_9_n671, mult_9_n669, mult_9_n676);
	and gate_mult_9_n665 (mult_9_n665, mult_9_n1054, mult_9_n1201);
	xor gate_mult_9_n666 (mult_9_n666, mult_9_n1201, mult_9_n1054);
	xor gate_mult_9_n662 (mult_9_n662, mult_9_n1153, mult_9_n1137);
	and gate_mult_9_n661 (mult_9_n661, mult_9_n1137, mult_9_n1153);
	and gate_mult_9_n660 (mult_9_n660, mult_9_n662, mult_9_n1121);
	or gate_mult_9_n663 (mult_9_n663, mult_9_n661, mult_9_n660);
	xor gate_mult_9_n664 (mult_9_n664, mult_9_n1121, mult_9_n662);
	xor gate_mult_9_n657 (mult_9_n657, mult_9_n1185, mult_9_n1169);
	and gate_mult_9_n656 (mult_9_n656, mult_9_n1169, mult_9_n1185);
	and gate_mult_9_n655 (mult_9_n655, mult_9_n666, mult_9_n657);
	or gate_mult_9_n658 (mult_9_n658, mult_9_n656, mult_9_n655);
	xor gate_mult_9_n659 (mult_9_n659, mult_9_n657, mult_9_n666);
	xor gate_mult_9_n652 (mult_9_n652, mult_9_n685, mult_9_n680);
	and gate_mult_9_n651 (mult_9_n651, mult_9_n680, mult_9_n685);
	and gate_mult_9_n650 (mult_9_n650, mult_9_n652, mult_9_n664);
	or gate_mult_9_n653 (mult_9_n653, mult_9_n651, mult_9_n650);
	xor gate_mult_9_n654 (mult_9_n654, mult_9_n664, mult_9_n652);
	xor gate_mult_9_n647 (mult_9_n647, mult_9_n659, mult_9_n675);
	and gate_mult_9_n646 (mult_9_n646, mult_9_n675, mult_9_n659);
	and gate_mult_9_n645 (mult_9_n645, mult_9_n647, mult_9_n654);
	or gate_mult_9_n648 (mult_9_n648, mult_9_n646, mult_9_n645);
	xor gate_mult_9_n649 (mult_9_n649, mult_9_n654, mult_9_n647);
	xor gate_mult_9_n642 (mult_9_n642, mult_9_n1200, mult_9_n1184);
	and gate_mult_9_n641 (mult_9_n641, mult_9_n1184, mult_9_n1200);
	and gate_mult_9_n640 (mult_9_n640, mult_9_n642, mult_9_n1168);
	or gate_mult_9_n643 (mult_9_n643, mult_9_n641, mult_9_n640);
	xor gate_mult_9_n644 (mult_9_n644, mult_9_n1168, mult_9_n642);
	xor gate_mult_9_n637 (mult_9_n637, mult_9_n1152, mult_9_n1136);
	and gate_mult_9_n636 (mult_9_n636, mult_9_n1136, mult_9_n1152);
	and gate_mult_9_n635 (mult_9_n635, mult_9_n637, mult_9_n1120);
	or gate_mult_9_n638 (mult_9_n638, mult_9_n636, mult_9_n635);
	xor gate_mult_9_n639 (mult_9_n639, mult_9_n1120, mult_9_n637);
	xor gate_mult_9_n632 (mult_9_n632, mult_9_n1104, mult_9_n665);
	and gate_mult_9_n631 (mult_9_n631, mult_9_n665, mult_9_n1104);
	and gate_mult_9_n630 (mult_9_n630, mult_9_n663, mult_9_n632);
	or gate_mult_9_n633 (mult_9_n633, mult_9_n631, mult_9_n630);
	xor gate_mult_9_n634 (mult_9_n634, mult_9_n632, mult_9_n663);
	xor gate_mult_9_n627 (mult_9_n627, mult_9_n658, mult_9_n644);
	and gate_mult_9_n626 (mult_9_n626, mult_9_n644, mult_9_n658);
	and gate_mult_9_n625 (mult_9_n625, mult_9_n627, mult_9_n639);
	or gate_mult_9_n628 (mult_9_n628, mult_9_n626, mult_9_n625);
	xor gate_mult_9_n629 (mult_9_n629, mult_9_n639, mult_9_n627);
	xor gate_mult_9_n622 (mult_9_n622, mult_9_n634, mult_9_n653);
	and gate_mult_9_n621 (mult_9_n621, mult_9_n653, mult_9_n634);
	and gate_mult_9_n620 (mult_9_n620, mult_9_n622, mult_9_n629);
	or gate_mult_9_n623 (mult_9_n623, mult_9_n621, mult_9_n620);
	xor gate_mult_9_n624 (mult_9_n624, mult_9_n629, mult_9_n622);
	and gate_mult_9_n618 (mult_9_n618, mult_9_n1053, mult_9_n1199);
	xor gate_mult_9_n619 (mult_9_n619, mult_9_n1199, mult_9_n1053);
	xor gate_mult_9_n615 (mult_9_n615, mult_9_n1135, mult_9_n1151);
	and gate_mult_9_n614 (mult_9_n614, mult_9_n1151, mult_9_n1135);
	and gate_mult_9_n613 (mult_9_n613, mult_9_n615, mult_9_n1119);
	or gate_mult_9_n616 (mult_9_n616, mult_9_n614, mult_9_n613);
	xor gate_mult_9_n617 (mult_9_n617, mult_9_n1119, mult_9_n615);
	xor gate_mult_9_n610 (mult_9_n610, mult_9_n1183, mult_9_n1167);
	and gate_mult_9_n609 (mult_9_n609, mult_9_n1167, mult_9_n1183);
	and gate_mult_9_n608 (mult_9_n608, mult_9_n610, mult_9_n1103);
	or gate_mult_9_n611 (mult_9_n611, mult_9_n609, mult_9_n608);
	xor gate_mult_9_n612 (mult_9_n612, mult_9_n1103, mult_9_n610);
	xor gate_mult_9_n605 (mult_9_n605, mult_9_n619, mult_9_n643);
	and gate_mult_9_n604 (mult_9_n604, mult_9_n643, mult_9_n619);
	and gate_mult_9_n603 (mult_9_n603, mult_9_n605, mult_9_n638);
	or gate_mult_9_n606 (mult_9_n606, mult_9_n604, mult_9_n603);
	xor gate_mult_9_n607 (mult_9_n607, mult_9_n638, mult_9_n605);
	xor gate_mult_9_n600 (mult_9_n600, mult_9_n612, mult_9_n617);
	and gate_mult_9_n599 (mult_9_n599, mult_9_n617, mult_9_n612);
	and gate_mult_9_n598 (mult_9_n598, mult_9_n600, mult_9_n633);
	or gate_mult_9_n601 (mult_9_n601, mult_9_n599, mult_9_n598);
	xor gate_mult_9_n602 (mult_9_n602, mult_9_n633, mult_9_n600);
	xor gate_mult_9_n595 (mult_9_n595, mult_9_n607, mult_9_n628);
	and gate_mult_9_n594 (mult_9_n594, mult_9_n628, mult_9_n607);
	and gate_mult_9_n593 (mult_9_n593, mult_9_n595, mult_9_n602);
	or gate_mult_9_n596 (mult_9_n596, mult_9_n594, mult_9_n593);
	xor gate_mult_9_n597 (mult_9_n597, mult_9_n602, mult_9_n595);
	xor gate_mult_9_n590 (mult_9_n590, mult_9_n1198, mult_9_n1182);
	and gate_mult_9_n589 (mult_9_n589, mult_9_n1182, mult_9_n1198);
	and gate_mult_9_n588 (mult_9_n588, mult_9_n590, mult_9_n1166);
	or gate_mult_9_n591 (mult_9_n591, mult_9_n589, mult_9_n588);
	xor gate_mult_9_n592 (mult_9_n592, mult_9_n1166, mult_9_n590);
	xor gate_mult_9_n585 (mult_9_n585, mult_9_n1150, mult_9_n1134);
	and gate_mult_9_n584 (mult_9_n584, mult_9_n1134, mult_9_n1150);
	and gate_mult_9_n583 (mult_9_n583, mult_9_n585, mult_9_n1118);
	or gate_mult_9_n586 (mult_9_n586, mult_9_n584, mult_9_n583);
	xor gate_mult_9_n587 (mult_9_n587, mult_9_n1118, mult_9_n585);
	xor gate_mult_9_n580 (mult_9_n580, mult_9_n1102, mult_9_n1086);
	and gate_mult_9_n579 (mult_9_n579, mult_9_n1086, mult_9_n1102);
	and gate_mult_9_n578 (mult_9_n578, mult_9_n580, mult_9_n618);
	or gate_mult_9_n581 (mult_9_n581, mult_9_n579, mult_9_n578);
	xor gate_mult_9_n582 (mult_9_n582, mult_9_n618, mult_9_n580);
	xor gate_mult_9_n575 (mult_9_n575, mult_9_n616, mult_9_n611);
	and gate_mult_9_n574 (mult_9_n574, mult_9_n611, mult_9_n616);
	and gate_mult_9_n573 (mult_9_n573, mult_9_n575, mult_9_n592);
	or gate_mult_9_n576 (mult_9_n576, mult_9_n574, mult_9_n573);
	xor gate_mult_9_n577 (mult_9_n577, mult_9_n592, mult_9_n575);
	xor gate_mult_9_n570 (mult_9_n570, mult_9_n587, mult_9_n582);
	and gate_mult_9_n569 (mult_9_n569, mult_9_n582, mult_9_n587);
	and gate_mult_9_n568 (mult_9_n568, mult_9_n606, mult_9_n570);
	or gate_mult_9_n571 (mult_9_n571, mult_9_n569, mult_9_n568);
	xor gate_mult_9_n572 (mult_9_n572, mult_9_n570, mult_9_n606);
	xor gate_mult_9_n565 (mult_9_n565, mult_9_n577, mult_9_n601);
	and gate_mult_9_n564 (mult_9_n564, mult_9_n601, mult_9_n577);
	and gate_mult_9_n563 (mult_9_n563, mult_9_n565, mult_9_n572);
	or gate_mult_9_n566 (mult_9_n566, mult_9_n564, mult_9_n563);
	xor gate_mult_9_n567 (mult_9_n567, mult_9_n572, mult_9_n565);
	and gate_mult_9_n561 (mult_9_n561, mult_9_n1052, mult_9_n1197);
	xor gate_mult_9_n562 (mult_9_n562, mult_9_n1197, mult_9_n1052);
	xor gate_mult_9_n558 (mult_9_n558, mult_9_n1133, mult_9_n1117);
	and gate_mult_9_n557 (mult_9_n557, mult_9_n1117, mult_9_n1133);
	and gate_mult_9_n556 (mult_9_n556, mult_9_n558, mult_9_n1101);
	or gate_mult_9_n559 (mult_9_n559, mult_9_n557, mult_9_n556);
	xor gate_mult_9_n560 (mult_9_n560, mult_9_n1101, mult_9_n558);
	xor gate_mult_9_n553 (mult_9_n553, mult_9_n1085, mult_9_n1149);
	and gate_mult_9_n552 (mult_9_n552, mult_9_n1149, mult_9_n1085);
	and gate_mult_9_n551 (mult_9_n551, mult_9_n553, mult_9_n1181);
	or gate_mult_9_n554 (mult_9_n554, mult_9_n552, mult_9_n551);
	xor gate_mult_9_n555 (mult_9_n555, mult_9_n1181, mult_9_n553);
	xor gate_mult_9_n548 (mult_9_n548, mult_9_n1165, mult_9_n562);
	and gate_mult_9_n547 (mult_9_n547, mult_9_n562, mult_9_n1165);
	and gate_mult_9_n546 (mult_9_n546, mult_9_n548, mult_9_n591);
	or gate_mult_9_n549 (mult_9_n549, mult_9_n547, mult_9_n546);
	xor gate_mult_9_n550 (mult_9_n550, mult_9_n591, mult_9_n548);
	xor gate_mult_9_n543 (mult_9_n543, mult_9_n586, mult_9_n581);
	and gate_mult_9_n542 (mult_9_n542, mult_9_n581, mult_9_n586);
	and gate_mult_9_n541 (mult_9_n541, mult_9_n543, mult_9_n555);
	or gate_mult_9_n544 (mult_9_n544, mult_9_n542, mult_9_n541);
	xor gate_mult_9_n545 (mult_9_n545, mult_9_n555, mult_9_n543);
	xor gate_mult_9_n538 (mult_9_n538, mult_9_n560, mult_9_n550);
	and gate_mult_9_n537 (mult_9_n537, mult_9_n550, mult_9_n560);
	and gate_mult_9_n536 (mult_9_n536, mult_9_n538, mult_9_n576);
	or gate_mult_9_n539 (mult_9_n539, mult_9_n537, mult_9_n536);
	xor gate_mult_9_n540 (mult_9_n540, mult_9_n576, mult_9_n538);
	xor gate_mult_9_n533 (mult_9_n533, mult_9_n545, mult_9_n571);
	and gate_mult_9_n532 (mult_9_n532, mult_9_n571, mult_9_n545);
	and gate_mult_9_n531 (mult_9_n531, mult_9_n540, mult_9_n533);
	or gate_mult_9_n534 (mult_9_n534, mult_9_n532, mult_9_n531);
	xor gate_mult_9_n535 (mult_9_n535, mult_9_n533, mult_9_n540);
	xor gate_mult_9_n528 (mult_9_n528, mult_9_n1068, mult_9_n1196);
	and gate_mult_9_n527 (mult_9_n527, mult_9_n1196, mult_9_n1068);
	and gate_mult_9_n526 (mult_9_n526, mult_9_n528, mult_9_n1180);
	or gate_mult_9_n529 (mult_9_n529, mult_9_n527, mult_9_n526);
	xor gate_mult_9_n530 (mult_9_n530, mult_9_n1180, mult_9_n528);
	xor gate_mult_9_n523 (mult_9_n523, mult_9_n1164, mult_9_n1148);
	and gate_mult_9_n522 (mult_9_n522, mult_9_n1148, mult_9_n1164);
	and gate_mult_9_n521 (mult_9_n521, mult_9_n523, mult_9_n1132);
	or gate_mult_9_n524 (mult_9_n524, mult_9_n522, mult_9_n521);
	xor gate_mult_9_n525 (mult_9_n525, mult_9_n1132, mult_9_n523);
	xor gate_mult_9_n518 (mult_9_n518, mult_9_n1116, mult_9_n1100);
	and gate_mult_9_n517 (mult_9_n517, mult_9_n1100, mult_9_n1116);
	and gate_mult_9_n516 (mult_9_n516, mult_9_n518, mult_9_n1084);
	or gate_mult_9_n519 (mult_9_n519, mult_9_n517, mult_9_n516);
	xor gate_mult_9_n520 (mult_9_n520, mult_9_n1084, mult_9_n518);
	xor gate_mult_9_n513 (mult_9_n513, mult_9_n561, mult_9_n559);
	and gate_mult_9_n512 (mult_9_n512, mult_9_n559, mult_9_n561);
	and gate_mult_9_n511 (mult_9_n511, mult_9_n513, mult_9_n554);
	or gate_mult_9_n514 (mult_9_n514, mult_9_n512, mult_9_n511);
	xor gate_mult_9_n515 (mult_9_n515, mult_9_n554, mult_9_n513);
	xor gate_mult_9_n508 (mult_9_n508, mult_9_n530, mult_9_n520);
	and gate_mult_9_n507 (mult_9_n507, mult_9_n520, mult_9_n530);
	and gate_mult_9_n506 (mult_9_n506, mult_9_n508, mult_9_n525);
	or gate_mult_9_n509 (mult_9_n509, mult_9_n507, mult_9_n506);
	xor gate_mult_9_n510 (mult_9_n510, mult_9_n525, mult_9_n508);
	xor gate_mult_9_n503 (mult_9_n503, mult_9_n549, mult_9_n544);
	and gate_mult_9_n502 (mult_9_n502, mult_9_n544, mult_9_n549);
	and gate_mult_9_n501 (mult_9_n501, mult_9_n503, mult_9_n515);
	or gate_mult_9_n504 (mult_9_n504, mult_9_n502, mult_9_n501);
	xor gate_mult_9_n505 (mult_9_n505, mult_9_n515, mult_9_n503);
	xor gate_mult_9_n498 (mult_9_n498, mult_9_n510, mult_9_n539);
	and gate_mult_9_n497 (mult_9_n497, mult_9_n539, mult_9_n510);
	and gate_mult_9_n496 (mult_9_n496, mult_9_n498, mult_9_n505);
	or gate_mult_9_n499 (mult_9_n499, mult_9_n497, mult_9_n496);
	xor gate_mult_9_n500 (mult_9_n500, mult_9_n505, mult_9_n498);
	not gate_mult_9_n495 (mult_9_n495, mult_9_n458);
	xor gate_mult_9_n492 (mult_9_n492, mult_9_n495, mult_9_n1099);
	and gate_mult_9_n491 (mult_9_n491, mult_9_n1099, mult_9_n495);
	and gate_mult_9_n490 (mult_9_n490, mult_9_n492, mult_9_n1147);
	or gate_mult_9_n493 (mult_9_n493, mult_9_n491, mult_9_n490);
	xor gate_mult_9_n494 (mult_9_n494, mult_9_n1147, mult_9_n492);
	xor gate_mult_9_n487 (mult_9_n487, mult_9_n1131, mult_9_n1163);
	and gate_mult_9_n486 (mult_9_n486, mult_9_n1163, mult_9_n1131);
	and gate_mult_9_n485 (mult_9_n485, mult_9_n487, mult_9_n1115);
	or gate_mult_9_n488 (mult_9_n488, mult_9_n486, mult_9_n485);
	xor gate_mult_9_n489 (mult_9_n489, mult_9_n1115, mult_9_n487);
	xor gate_mult_9_n482 (mult_9_n482, mult_9_n1179, mult_9_n1083);
	and gate_mult_9_n481 (mult_9_n481, mult_9_n1083, mult_9_n1179);
	and gate_mult_9_n480 (mult_9_n480, mult_9_n482, mult_9_n1195);
	or gate_mult_9_n483 (mult_9_n483, mult_9_n481, mult_9_n480);
	xor gate_mult_9_n484 (mult_9_n484, mult_9_n1195, mult_9_n482);
	xor gate_mult_9_n477 (mult_9_n477, mult_9_n529, mult_9_n524);
	and gate_mult_9_n476 (mult_9_n476, mult_9_n524, mult_9_n529);
	and gate_mult_9_n475 (mult_9_n475, mult_9_n477, mult_9_n519);
	or gate_mult_9_n478 (mult_9_n478, mult_9_n476, mult_9_n475);
	xor gate_mult_9_n479 (mult_9_n479, mult_9_n519, mult_9_n477);
	xor gate_mult_9_n472 (mult_9_n472, mult_9_n494, mult_9_n484);
	and gate_mult_9_n471 (mult_9_n471, mult_9_n484, mult_9_n494);
	and gate_mult_9_n470 (mult_9_n470, mult_9_n472, mult_9_n489);
	or gate_mult_9_n473 (mult_9_n473, mult_9_n471, mult_9_n470);
	xor gate_mult_9_n474 (mult_9_n474, mult_9_n489, mult_9_n472);
	xor gate_mult_9_n467 (mult_9_n467, mult_9_n514, mult_9_n479);
	and gate_mult_9_n466 (mult_9_n466, mult_9_n479, mult_9_n514);
	and gate_mult_9_n465 (mult_9_n465, mult_9_n467, mult_9_n509);
	or gate_mult_9_n468 (mult_9_n468, mult_9_n466, mult_9_n465);
	xor gate_mult_9_n469 (mult_9_n469, mult_9_n509, mult_9_n467);
	xor gate_mult_9_n462 (mult_9_n462, mult_9_n474, mult_9_n504);
	and gate_mult_9_n461 (mult_9_n461, mult_9_n504, mult_9_n474);
	and gate_mult_9_n460 (mult_9_n460, mult_9_n462, mult_9_n469);
	or gate_mult_9_n463 (mult_9_n463, mult_9_n461, mult_9_n460);
	xor gate_mult_9_n464 (mult_9_n464, mult_9_n469, mult_9_n462);
	not gate_mult_9_n459 (mult_9_n459, mult_9_n458);
	xor gate_mult_9_n455 (mult_9_n455, mult_9_n1067, mult_9_n459);
	and gate_mult_9_n454 (mult_9_n454, mult_9_n459, mult_9_n1067);
	and gate_mult_9_n453 (mult_9_n453, mult_9_n455, mult_9_n1178);
	or gate_mult_9_n456 (mult_9_n456, mult_9_n454, mult_9_n453);
	xor gate_mult_9_n457 (mult_9_n457, mult_9_n1178, mult_9_n455);
	xor gate_mult_9_n450 (mult_9_n450, mult_9_n1114, mult_9_n1098);
	and gate_mult_9_n449 (mult_9_n449, mult_9_n1098, mult_9_n1114);
	and gate_mult_9_n448 (mult_9_n448, mult_9_n450, mult_9_n1130);
	or gate_mult_9_n451 (mult_9_n451, mult_9_n449, mult_9_n448);
	xor gate_mult_9_n452 (mult_9_n452, mult_9_n1130, mult_9_n450);
	xor gate_mult_9_n445 (mult_9_n445, mult_9_n1162, mult_9_n1146);
	and gate_mult_9_n444 (mult_9_n444, mult_9_n1146, mult_9_n1162);
	and gate_mult_9_n443 (mult_9_n443, mult_9_n445, mult_9_n1082);
	or gate_mult_9_n446 (mult_9_n446, mult_9_n444, mult_9_n443);
	xor gate_mult_9_n447 (mult_9_n447, mult_9_n1082, mult_9_n445);
	xor gate_mult_9_n440 (mult_9_n440, mult_9_n457, mult_9_n493);
	and gate_mult_9_n439 (mult_9_n439, mult_9_n493, mult_9_n457);
	and gate_mult_9_n438 (mult_9_n438, mult_9_n440, mult_9_n488);
	or gate_mult_9_n441 (mult_9_n441, mult_9_n439, mult_9_n438);
	xor gate_mult_9_n442 (mult_9_n442, mult_9_n488, mult_9_n440);
	xor gate_mult_9_n435 (mult_9_n435, mult_9_n483, mult_9_n447);
	and gate_mult_9_n434 (mult_9_n434, mult_9_n447, mult_9_n483);
	and gate_mult_9_n433 (mult_9_n433, mult_9_n435, mult_9_n452);
	or gate_mult_9_n436 (mult_9_n436, mult_9_n434, mult_9_n433);
	xor gate_mult_9_n437 (mult_9_n437, mult_9_n452, mult_9_n435);
	xor gate_mult_9_n430 (mult_9_n430, mult_9_n478, mult_9_n442);
	and gate_mult_9_n429 (mult_9_n429, mult_9_n442, mult_9_n478);
	and gate_mult_9_n428 (mult_9_n428, mult_9_n430, mult_9_n473);
	or gate_mult_9_n431 (mult_9_n431, mult_9_n429, mult_9_n428);
	xor gate_mult_9_n432 (mult_9_n432, mult_9_n473, mult_9_n430);
	xor gate_mult_9_n425 (mult_9_n425, mult_9_n437, mult_9_n468);
	and gate_mult_9_n424 (mult_9_n424, mult_9_n468, mult_9_n437);
	and gate_mult_9_n423 (mult_9_n423, mult_9_n425, mult_9_n432);
	or gate_mult_9_n426 (mult_9_n426, mult_9_n424, mult_9_n423);
	xor gate_mult_9_n427 (mult_9_n427, mult_9_n432, mult_9_n425);
	xor gate_mult_9_n420 (mult_9_n420, mult_9_n458, mult_9_n1066);
	and gate_mult_9_n419 (mult_9_n419, mult_9_n1066, mult_9_n458);
	and gate_mult_9_n418 (mult_9_n418, mult_9_n420, mult_9_n1129);
	or gate_mult_9_n421 (mult_9_n421, mult_9_n419, mult_9_n418);
	xor gate_mult_9_n422 (mult_9_n422, mult_9_n1129, mult_9_n420);
	xor gate_mult_9_n415 (mult_9_n415, mult_9_n1113, mult_9_n1097);
	and gate_mult_9_n414 (mult_9_n414, mult_9_n1097, mult_9_n1113);
	and gate_mult_9_n413 (mult_9_n413, mult_9_n415, mult_9_n1145);
	or gate_mult_9_n416 (mult_9_n416, mult_9_n414, mult_9_n413);
	xor gate_mult_9_n417 (mult_9_n417, mult_9_n1145, mult_9_n415);
	xor gate_mult_9_n410 (mult_9_n410, mult_9_n1161, mult_9_n1081);
	and gate_mult_9_n409 (mult_9_n409, mult_9_n1081, mult_9_n1161);
	and gate_mult_9_n408 (mult_9_n408, mult_9_n410, mult_9_n1177);
	or gate_mult_9_n411 (mult_9_n411, mult_9_n409, mult_9_n408);
	xor gate_mult_9_n412 (mult_9_n412, mult_9_n1177, mult_9_n410);
	xor gate_mult_9_n405 (mult_9_n405, mult_9_n456, mult_9_n422);
	and gate_mult_9_n404 (mult_9_n404, mult_9_n422, mult_9_n456);
	and gate_mult_9_n403 (mult_9_n403, mult_9_n405, mult_9_n451);
	or gate_mult_9_n406 (mult_9_n406, mult_9_n404, mult_9_n403);
	xor gate_mult_9_n407 (mult_9_n407, mult_9_n451, mult_9_n405);
	xor gate_mult_9_n400 (mult_9_n400, mult_9_n446, mult_9_n412);
	and gate_mult_9_n399 (mult_9_n399, mult_9_n412, mult_9_n446);
	and gate_mult_9_n398 (mult_9_n398, mult_9_n400, mult_9_n417);
	or gate_mult_9_n401 (mult_9_n401, mult_9_n399, mult_9_n398);
	xor gate_mult_9_n402 (mult_9_n402, mult_9_n417, mult_9_n400);
	xor gate_mult_9_n395 (mult_9_n395, mult_9_n407, mult_9_n441);
	and gate_mult_9_n394 (mult_9_n394, mult_9_n441, mult_9_n407);
	and gate_mult_9_n393 (mult_9_n393, mult_9_n395, mult_9_n436);
	or gate_mult_9_n396 (mult_9_n396, mult_9_n394, mult_9_n393);
	xor gate_mult_9_n397 (mult_9_n397, mult_9_n436, mult_9_n395);
	xor gate_mult_9_n390 (mult_9_n390, mult_9_n402, mult_9_n431);
	and gate_mult_9_n389 (mult_9_n389, mult_9_n431, mult_9_n402);
	and gate_mult_9_n388 (mult_9_n388, mult_9_n390, mult_9_n397);
	or gate_mult_9_n391 (mult_9_n391, mult_9_n389, mult_9_n388);
	xor gate_mult_9_n392 (mult_9_n392, mult_9_n397, mult_9_n390);
	not gate_mult_9_n387 (mult_9_n387, mult_9_n386);
	xor gate_mult_9_n383 (mult_9_n383, mult_9_n387, mult_9_n1160);
	and gate_mult_9_n382 (mult_9_n382, mult_9_n1160, mult_9_n387);
	and gate_mult_9_n381 (mult_9_n381, mult_9_n383, mult_9_n1144);
	or gate_mult_9_n384 (mult_9_n384, mult_9_n382, mult_9_n381);
	xor gate_mult_9_n385 (mult_9_n385, mult_9_n1144, mult_9_n383);
	xor gate_mult_9_n378 (mult_9_n378, mult_9_n1128, mult_9_n1112);
	and gate_mult_9_n377 (mult_9_n377, mult_9_n1112, mult_9_n1128);
	and gate_mult_9_n376 (mult_9_n376, mult_9_n378, mult_9_n1080);
	or gate_mult_9_n379 (mult_9_n379, mult_9_n377, mult_9_n376);
	xor gate_mult_9_n380 (mult_9_n380, mult_9_n1080, mult_9_n378);
	xor gate_mult_9_n373 (mult_9_n373, mult_9_n1096, mult_9_n421);
	and gate_mult_9_n372 (mult_9_n372, mult_9_n421, mult_9_n1096);
	and gate_mult_9_n371 (mult_9_n371, mult_9_n416, mult_9_n373);
	or gate_mult_9_n374 (mult_9_n374, mult_9_n372, mult_9_n371);
	xor gate_mult_9_n375 (mult_9_n375, mult_9_n373, mult_9_n416);
	xor gate_mult_9_n368 (mult_9_n368, mult_9_n411, mult_9_n385);
	and gate_mult_9_n367 (mult_9_n367, mult_9_n385, mult_9_n411);
	and gate_mult_9_n366 (mult_9_n366, mult_9_n368, mult_9_n380);
	or gate_mult_9_n369 (mult_9_n369, mult_9_n367, mult_9_n366);
	xor gate_mult_9_n370 (mult_9_n370, mult_9_n380, mult_9_n368);
	xor gate_mult_9_n363 (mult_9_n363, mult_9_n375, mult_9_n406);
	and gate_mult_9_n362 (mult_9_n362, mult_9_n406, mult_9_n375);
	and gate_mult_9_n361 (mult_9_n361, mult_9_n363, mult_9_n401);
	or gate_mult_9_n364 (mult_9_n364, mult_9_n362, mult_9_n361);
	xor gate_mult_9_n365 (mult_9_n365, mult_9_n401, mult_9_n363);
	xor gate_mult_9_n358 (mult_9_n358, mult_9_n370, mult_9_n365);
	and gate_mult_9_n357 (mult_9_n357, mult_9_n365, mult_9_n370);
	and gate_mult_9_n356 (mult_9_n356, mult_9_n358, mult_9_n396);
	or gate_mult_9_n359 (mult_9_n359, mult_9_n357, mult_9_n356);
	xor gate_mult_9_n360 (mult_9_n360, mult_9_n396, mult_9_n358);
	xor gate_mult_9_n353 (mult_9_n353, mult_9_n386, mult_9_n1065);
	and gate_mult_9_n352 (mult_9_n352, mult_9_n1065, mult_9_n386);
	and gate_mult_9_n351 (mult_9_n351, mult_9_n353, mult_9_n1127);
	or gate_mult_9_n354 (mult_9_n354, mult_9_n352, mult_9_n351);
	xor gate_mult_9_n355 (mult_9_n355, mult_9_n1127, mult_9_n353);
	xor gate_mult_9_n348 (mult_9_n348, mult_9_n1095, mult_9_n1111);
	and gate_mult_9_n347 (mult_9_n347, mult_9_n1111, mult_9_n1095);
	and gate_mult_9_n346 (mult_9_n346, mult_9_n348, mult_9_n1079);
	or gate_mult_9_n349 (mult_9_n349, mult_9_n347, mult_9_n346);
	xor gate_mult_9_n350 (mult_9_n350, mult_9_n1079, mult_9_n348);
	xor gate_mult_9_n343 (mult_9_n343, mult_9_n1143, mult_9_n1159);
	and gate_mult_9_n342 (mult_9_n342, mult_9_n1159, mult_9_n1143);
	and gate_mult_9_n341 (mult_9_n341, mult_9_n355, mult_9_n343);
	or gate_mult_9_n344 (mult_9_n344, mult_9_n342, mult_9_n341);
	xor gate_mult_9_n345 (mult_9_n345, mult_9_n343, mult_9_n355);
	xor gate_mult_9_n338 (mult_9_n338, mult_9_n384, mult_9_n379);
	and gate_mult_9_n337 (mult_9_n337, mult_9_n379, mult_9_n384);
	and gate_mult_9_n336 (mult_9_n336, mult_9_n338, mult_9_n350);
	or gate_mult_9_n339 (mult_9_n339, mult_9_n337, mult_9_n336);
	xor gate_mult_9_n340 (mult_9_n340, mult_9_n350, mult_9_n338);
	xor gate_mult_9_n333 (mult_9_n333, mult_9_n345, mult_9_n374);
	and gate_mult_9_n332 (mult_9_n332, mult_9_n374, mult_9_n345);
	and gate_mult_9_n331 (mult_9_n331, mult_9_n369, mult_9_n333);
	or gate_mult_9_n334 (mult_9_n334, mult_9_n332, mult_9_n331);
	xor gate_mult_9_n335 (mult_9_n335, mult_9_n333, mult_9_n369);
	xor gate_mult_9_n328 (mult_9_n328, mult_9_n340, mult_9_n364);
	and gate_mult_9_n327 (mult_9_n327, mult_9_n364, mult_9_n340);
	and gate_mult_9_n326 (mult_9_n326, mult_9_n328, mult_9_n335);
	or gate_mult_9_n329 (mult_9_n329, mult_9_n327, mult_9_n326);
	xor gate_mult_9_n330 (mult_9_n330, mult_9_n335, mult_9_n328);
	not gate_mult_9_n325 (mult_9_n325, mult_9_n324);
	xor gate_mult_9_n321 (mult_9_n321, mult_9_n325, mult_9_n1142);
	and gate_mult_9_n320 (mult_9_n320, mult_9_n1142, mult_9_n325);
	and gate_mult_9_n319 (mult_9_n319, mult_9_n321, mult_9_n1126);
	or gate_mult_9_n322 (mult_9_n322, mult_9_n320, mult_9_n319);
	xor gate_mult_9_n323 (mult_9_n323, mult_9_n1126, mult_9_n321);
	xor gate_mult_9_n316 (mult_9_n316, mult_9_n1110, mult_9_n1094);
	and gate_mult_9_n315 (mult_9_n315, mult_9_n1094, mult_9_n1110);
	and gate_mult_9_n314 (mult_9_n314, mult_9_n316, mult_9_n1078);
	or gate_mult_9_n317 (mult_9_n317, mult_9_n315, mult_9_n314);
	xor gate_mult_9_n318 (mult_9_n318, mult_9_n1078, mult_9_n316);
	xor gate_mult_9_n311 (mult_9_n311, mult_9_n354, mult_9_n349);
	and gate_mult_9_n310 (mult_9_n310, mult_9_n349, mult_9_n354);
	and gate_mult_9_n309 (mult_9_n309, mult_9_n311, mult_9_n344);
	or gate_mult_9_n312 (mult_9_n312, mult_9_n310, mult_9_n309);
	xor gate_mult_9_n313 (mult_9_n313, mult_9_n344, mult_9_n311);
	xor gate_mult_9_n306 (mult_9_n306, mult_9_n323, mult_9_n318);
	and gate_mult_9_n305 (mult_9_n305, mult_9_n318, mult_9_n323);
	and gate_mult_9_n304 (mult_9_n304, mult_9_n339, mult_9_n306);
	or gate_mult_9_n307 (mult_9_n307, mult_9_n305, mult_9_n304);
	xor gate_mult_9_n308 (mult_9_n308, mult_9_n306, mult_9_n339);
	xor gate_mult_9_n301 (mult_9_n301, mult_9_n313, mult_9_n334);
	and gate_mult_9_n300 (mult_9_n300, mult_9_n334, mult_9_n313);
	and gate_mult_9_n299 (mult_9_n299, mult_9_n301, mult_9_n308);
	or gate_mult_9_n302 (mult_9_n302, mult_9_n300, mult_9_n299);
	xor gate_mult_9_n303 (mult_9_n303, mult_9_n308, mult_9_n301);
	xor gate_mult_9_n296 (mult_9_n296, mult_9_n324, mult_9_n1064);
	and gate_mult_9_n295 (mult_9_n295, mult_9_n1064, mult_9_n324);
	and gate_mult_9_n294 (mult_9_n294, mult_9_n296, mult_9_n1109);
	or gate_mult_9_n297 (mult_9_n297, mult_9_n295, mult_9_n294);
	xor gate_mult_9_n298 (mult_9_n298, mult_9_n1109, mult_9_n296);
	xor gate_mult_9_n291 (mult_9_n291, mult_9_n1093, mult_9_n1077);
	and gate_mult_9_n290 (mult_9_n290, mult_9_n1077, mult_9_n1093);
	and gate_mult_9_n289 (mult_9_n289, mult_9_n291, mult_9_n1125);
	or gate_mult_9_n292 (mult_9_n292, mult_9_n290, mult_9_n289);
	xor gate_mult_9_n293 (mult_9_n293, mult_9_n1125, mult_9_n291);
	xor gate_mult_9_n286 (mult_9_n286, mult_9_n1141, mult_9_n298);
	and gate_mult_9_n285 (mult_9_n285, mult_9_n298, mult_9_n1141);
	and gate_mult_9_n284 (mult_9_n284, mult_9_n286, mult_9_n322);
	or gate_mult_9_n287 (mult_9_n287, mult_9_n285, mult_9_n284);
	xor gate_mult_9_n288 (mult_9_n288, mult_9_n322, mult_9_n286);
	xor gate_mult_9_n281 (mult_9_n281, mult_9_n317, mult_9_n293);
	and gate_mult_9_n280 (mult_9_n280, mult_9_n293, mult_9_n317);
	and gate_mult_9_n279 (mult_9_n279, mult_9_n288, mult_9_n281);
	or gate_mult_9_n282 (mult_9_n282, mult_9_n280, mult_9_n279);
	xor gate_mult_9_n283 (mult_9_n283, mult_9_n281, mult_9_n288);
	xor gate_mult_9_n276 (mult_9_n276, mult_9_n312, mult_9_n307);
	and gate_mult_9_n275 (mult_9_n275, mult_9_n307, mult_9_n312);
	and gate_mult_9_n274 (mult_9_n274, mult_9_n276, mult_9_n283);
	or gate_mult_9_n277 (mult_9_n277, mult_9_n275, mult_9_n274);
	xor gate_mult_9_n278 (mult_9_n278, mult_9_n283, mult_9_n276);
	not gate_mult_9_n273 (mult_9_n273, mult_9_n272);
	xor gate_mult_9_n269 (mult_9_n269, mult_9_n273, mult_9_n1124);
	and gate_mult_9_n268 (mult_9_n268, mult_9_n1124, mult_9_n273);
	and gate_mult_9_n267 (mult_9_n267, mult_9_n269, mult_9_n1108);
	or gate_mult_9_n270 (mult_9_n270, mult_9_n268, mult_9_n267);
	xor gate_mult_9_n271 (mult_9_n271, mult_9_n1108, mult_9_n269);
	xor gate_mult_9_n264 (mult_9_n264, mult_9_n1092, mult_9_n1076);
	and gate_mult_9_n263 (mult_9_n263, mult_9_n1076, mult_9_n1092);
	and gate_mult_9_n262 (mult_9_n262, mult_9_n264, mult_9_n297);
	or gate_mult_9_n265 (mult_9_n265, mult_9_n263, mult_9_n262);
	xor gate_mult_9_n266 (mult_9_n266, mult_9_n297, mult_9_n264);
	xor gate_mult_9_n259 (mult_9_n259, mult_9_n292, mult_9_n271);
	and gate_mult_9_n258 (mult_9_n258, mult_9_n271, mult_9_n292);
	and gate_mult_9_n257 (mult_9_n257, mult_9_n259, mult_9_n266);
	or gate_mult_9_n260 (mult_9_n260, mult_9_n258, mult_9_n257);
	xor gate_mult_9_n261 (mult_9_n261, mult_9_n266, mult_9_n259);
	xor gate_mult_9_n254 (mult_9_n254, mult_9_n287, mult_9_n282);
	and gate_mult_9_n253 (mult_9_n253, mult_9_n282, mult_9_n287);
	and gate_mult_9_n252 (mult_9_n252, mult_9_n254, mult_9_n261);
	or gate_mult_9_n255 (mult_9_n255, mult_9_n253, mult_9_n252);
	xor gate_mult_9_n256 (mult_9_n256, mult_9_n261, mult_9_n254);
	xor gate_mult_9_n249 (mult_9_n249, mult_9_n272, mult_9_n1063);
	and gate_mult_9_n248 (mult_9_n248, mult_9_n1063, mult_9_n272);
	and gate_mult_9_n247 (mult_9_n247, mult_9_n249, mult_9_n1107);
	or gate_mult_9_n250 (mult_9_n250, mult_9_n248, mult_9_n247);
	xor gate_mult_9_n251 (mult_9_n251, mult_9_n1107, mult_9_n249);
	xor gate_mult_9_n244 (mult_9_n244, mult_9_n1075, mult_9_n1091);
	and gate_mult_9_n243 (mult_9_n243, mult_9_n1091, mult_9_n1075);
	and gate_mult_9_n242 (mult_9_n242, mult_9_n244, mult_9_n1123);
	or gate_mult_9_n245 (mult_9_n245, mult_9_n243, mult_9_n242);
	xor gate_mult_9_n246 (mult_9_n246, mult_9_n1123, mult_9_n244);
	xor gate_mult_9_n239 (mult_9_n239, mult_9_n251, mult_9_n270);
	and gate_mult_9_n238 (mult_9_n238, mult_9_n270, mult_9_n251);
	and gate_mult_9_n237 (mult_9_n237, mult_9_n239, mult_9_n265);
	or gate_mult_9_n240 (mult_9_n240, mult_9_n238, mult_9_n237);
	xor gate_mult_9_n241 (mult_9_n241, mult_9_n265, mult_9_n239);
	xor gate_mult_9_n234 (mult_9_n234, mult_9_n246, mult_9_n241);
	and gate_mult_9_n233 (mult_9_n233, mult_9_n241, mult_9_n246);
	and gate_mult_9_n232 (mult_9_n232, mult_9_n234, mult_9_n260);
	or gate_mult_9_n235 (mult_9_n235, mult_9_n233, mult_9_n232);
	xor gate_mult_9_n236 (mult_9_n236, mult_9_n260, mult_9_n234);
	not gate_mult_9_n231 (mult_9_n231, mult_9_n230);
	xor gate_mult_9_n227 (mult_9_n227, mult_9_n231, mult_9_n1106);
	and gate_mult_9_n226 (mult_9_n226, mult_9_n1106, mult_9_n231);
	and gate_mult_9_n225 (mult_9_n225, mult_9_n227, mult_9_n1090);
	or gate_mult_9_n228 (mult_9_n228, mult_9_n226, mult_9_n225);
	xor gate_mult_9_n229 (mult_9_n229, mult_9_n1090, mult_9_n227);
	xor gate_mult_9_n222 (mult_9_n222, mult_9_n1074, mult_9_n250);
	and gate_mult_9_n221 (mult_9_n221, mult_9_n250, mult_9_n1074);
	and gate_mult_9_n220 (mult_9_n220, mult_9_n245, mult_9_n222);
	or gate_mult_9_n223 (mult_9_n223, mult_9_n221, mult_9_n220);
	xor gate_mult_9_n224 (mult_9_n224, mult_9_n222, mult_9_n245);
	xor gate_mult_9_n217 (mult_9_n217, mult_9_n229, mult_9_n224);
	and gate_mult_9_n216 (mult_9_n216, mult_9_n224, mult_9_n229);
	and gate_mult_9_n215 (mult_9_n215, mult_9_n217, mult_9_n240);
	or gate_mult_9_n218 (mult_9_n218, mult_9_n216, mult_9_n215);
	xor gate_mult_9_n219 (mult_9_n219, mult_9_n240, mult_9_n217);
	xor gate_mult_9_n212 (mult_9_n212, mult_9_n230, mult_9_n1062);
	and gate_mult_9_n211 (mult_9_n211, mult_9_n1062, mult_9_n230);
	and gate_mult_9_n210 (mult_9_n210, mult_9_n212, mult_9_n1089);
	or gate_mult_9_n213 (mult_9_n213, mult_9_n211, mult_9_n210);
	xor gate_mult_9_n214 (mult_9_n214, mult_9_n1089, mult_9_n212);
	xor gate_mult_9_n207 (mult_9_n207, mult_9_n1073, mult_9_n1105);
	and gate_mult_9_n206 (mult_9_n206, mult_9_n1105, mult_9_n1073);
	and gate_mult_9_n205 (mult_9_n205, mult_9_n214, mult_9_n207);
	or gate_mult_9_n208 (mult_9_n208, mult_9_n206, mult_9_n205);
	xor gate_mult_9_n209 (mult_9_n209, mult_9_n207, mult_9_n214);
	xor gate_mult_9_n202 (mult_9_n202, mult_9_n228, mult_9_n209);
	and gate_mult_9_n201 (mult_9_n201, mult_9_n209, mult_9_n228);
	and gate_mult_9_n200 (mult_9_n200, mult_9_n202, mult_9_n223);
	or gate_mult_9_n203 (mult_9_n203, mult_9_n201, mult_9_n200);
	xor gate_mult_9_n204 (mult_9_n204, mult_9_n223, mult_9_n202);
	not gate_mult_9_n199 (mult_9_n199, mult_9_n198);
	xor gate_mult_9_n195 (mult_9_n195, mult_9_n199, mult_9_n1088);
	and gate_mult_9_n194 (mult_9_n194, mult_9_n1088, mult_9_n199);
	and gate_mult_9_n193 (mult_9_n193, mult_9_n195, mult_9_n1072);
	or gate_mult_9_n196 (mult_9_n196, mult_9_n194, mult_9_n193);
	xor gate_mult_9_n197 (mult_9_n197, mult_9_n1072, mult_9_n195);
	xor gate_mult_9_n190 (mult_9_n190, mult_9_n213, mult_9_n208);
	and gate_mult_9_n189 (mult_9_n189, mult_9_n208, mult_9_n213);
	and gate_mult_9_n188 (mult_9_n188, mult_9_n190, mult_9_n197);
	or gate_mult_9_n191 (mult_9_n191, mult_9_n189, mult_9_n188);
	xor gate_mult_9_n192 (mult_9_n192, mult_9_n197, mult_9_n190);
	xor gate_mult_9_n185 (mult_9_n185, mult_9_n198, mult_9_n1061);
	and gate_mult_9_n184 (mult_9_n184, mult_9_n1061, mult_9_n198);
	and gate_mult_9_n183 (mult_9_n183, mult_9_n185, mult_9_n1071);
	or gate_mult_9_n186 (mult_9_n186, mult_9_n184, mult_9_n183);
	xor gate_mult_9_n187 (mult_9_n187, mult_9_n1071, mult_9_n185);
	xor gate_mult_9_n180 (mult_9_n180, mult_9_n1087, mult_9_n187);
	and gate_mult_9_n179 (mult_9_n179, mult_9_n187, mult_9_n1087);
	and gate_mult_9_n178 (mult_9_n178, mult_9_n180, mult_9_n196);
	or gate_mult_9_n181 (mult_9_n181, mult_9_n179, mult_9_n178);
	xor gate_mult_9_n182 (mult_9_n182, mult_9_n196, mult_9_n180);
	not gate_mult_9_n177 (mult_9_n177, mult_9_n176);
	xor gate_mult_9_n173 (mult_9_n173, mult_9_n177, mult_9_n1070);
	and gate_mult_9_n172 (mult_9_n172, mult_9_n1070, mult_9_n177);
	and gate_mult_9_n171 (mult_9_n171, mult_9_n173, mult_9_n186);
	or gate_mult_9_n174 (mult_9_n174, mult_9_n172, mult_9_n171);
	xor gate_mult_9_n175 (mult_9_n175, mult_9_n186, mult_9_n173);
	xor gate_mult_9_n169 (mult_9_n169, mult_9_n1069, mult_9_n1060);
	xor gate_mult_9_n170 (mult_9_n170, mult_9_n176, mult_9_n169);
	and gate_mult_9_n168 (mult_9_n168, mult_9_n1211, mult_9_n1059);
	xor gate_sum_1 (sum_1, mult_9_n1059, mult_9_n1211);
	xor gate_mult_9_n138 (mult_9_n138, mult_9_n1210, mult_9_n1194);
	and gate_mult_9_n137 (mult_9_n137, mult_9_n1194, mult_9_n1210);
	and gate_mult_9_n136 (mult_9_n136, mult_9_n138, mult_9_n168);
	or gate_mult_9_n167 (mult_9_n167, mult_9_n137, mult_9_n136);
	xor gate_sum_2 (sum_2, mult_9_n168, mult_9_n138);
	xor gate_mult_9_n135 (mult_9_n135, mult_9_n1058, mult_9_n754);
	and gate_mult_9_n134 (mult_9_n134, mult_9_n754, mult_9_n1058);
	and gate_mult_9_n133 (mult_9_n133, mult_9_n135, mult_9_n167);
	or gate_mult_9_n166 (mult_9_n166, mult_9_n134, mult_9_n133);
	xor gate_sum_3 (sum_3, mult_9_n167, mult_9_n135);
	xor gate_mult_9_n132 (mult_9_n132, mult_9_n753, mult_9_n752);
	and gate_mult_9_n131 (mult_9_n131, mult_9_n752, mult_9_n753);
	and gate_mult_9_n130 (mult_9_n130, mult_9_n132, mult_9_n166);
	or gate_mult_9_n165 (mult_9_n165, mult_9_n131, mult_9_n130);
	xor gate_sum_4 (sum_4, mult_9_n166, mult_9_n132);
	xor gate_mult_9_n129 (mult_9_n129, mult_9_n751, mult_9_n745);
	and gate_mult_9_n128 (mult_9_n128, mult_9_n745, mult_9_n751);
	and gate_mult_9_n127 (mult_9_n127, mult_9_n165, mult_9_n129);
	or gate_mult_9_n164 (mult_9_n164, mult_9_n128, mult_9_n127);
	xor gate_sum_5 (sum_5, mult_9_n129, mult_9_n165);
	xor gate_mult_9_n126 (mult_9_n126, mult_9_n740, mult_9_n735);
	and gate_mult_9_n125 (mult_9_n125, mult_9_n735, mult_9_n740);
	and gate_mult_9_n124 (mult_9_n124, mult_9_n164, mult_9_n126);
	or gate_mult_9_n163 (mult_9_n163, mult_9_n125, mult_9_n124);
	xor gate_sum_6 (sum_6, mult_9_n126, mult_9_n164);
	xor gate_mult_9_n123 (mult_9_n123, mult_9_n734, mult_9_n723);
	and gate_mult_9_n122 (mult_9_n122, mult_9_n723, mult_9_n734);
	and gate_mult_9_n121 (mult_9_n121, mult_9_n163, mult_9_n123);
	or gate_mult_9_n162 (mult_9_n162, mult_9_n122, mult_9_n121);
	xor gate_sum_7 (sum_7, mult_9_n123, mult_9_n163);
	xor gate_mult_9_n120 (mult_9_n120, mult_9_n722, mult_9_n708);
	and gate_mult_9_n119 (mult_9_n119, mult_9_n708, mult_9_n722);
	and gate_mult_9_n118 (mult_9_n118, mult_9_n162, mult_9_n120);
	or gate_mult_9_n161 (mult_9_n161, mult_9_n119, mult_9_n118);
	xor gate_sum_8 (sum_8, mult_9_n120, mult_9_n162);
	xor gate_mult_9_n117 (mult_9_n117, mult_9_n707, mult_9_n691);
	and gate_mult_9_n116 (mult_9_n116, mult_9_n691, mult_9_n707);
	and gate_mult_9_n115 (mult_9_n115, mult_9_n161, mult_9_n117);
	or gate_mult_9_n160 (mult_9_n160, mult_9_n116, mult_9_n115);
	xor gate_sum_9 (sum_9, mult_9_n117, mult_9_n161);
	xor gate_mult_9_n114 (mult_9_n114, mult_9_n690, mult_9_n671);
	and gate_mult_9_n113 (mult_9_n113, mult_9_n671, mult_9_n690);
	and gate_mult_9_n112 (mult_9_n112, mult_9_n160, mult_9_n114);
	or gate_mult_9_n159 (mult_9_n159, mult_9_n113, mult_9_n112);
	xor gate_sum_10 (sum_10, mult_9_n114, mult_9_n160);
	xor gate_mult_9_n111 (mult_9_n111, mult_9_n670, mult_9_n649);
	and gate_mult_9_n110 (mult_9_n110, mult_9_n649, mult_9_n670);
	and gate_mult_9_n109 (mult_9_n109, mult_9_n159, mult_9_n111);
	or gate_mult_9_n158 (mult_9_n158, mult_9_n110, mult_9_n109);
	xor gate_sum_11 (sum_11, mult_9_n111, mult_9_n159);
	xor gate_mult_9_n108 (mult_9_n108, mult_9_n648, mult_9_n624);
	and gate_mult_9_n107 (mult_9_n107, mult_9_n624, mult_9_n648);
	and gate_mult_9_n106 (mult_9_n106, mult_9_n158, mult_9_n108);
	or gate_mult_9_n157 (mult_9_n157, mult_9_n107, mult_9_n106);
	xor gate_sum_12 (sum_12, mult_9_n108, mult_9_n158);
	xor gate_mult_9_n105 (mult_9_n105, mult_9_n623, mult_9_n597);
	and gate_mult_9_n104 (mult_9_n104, mult_9_n597, mult_9_n623);
	and gate_mult_9_n103 (mult_9_n103, mult_9_n157, mult_9_n105);
	or gate_mult_9_n156 (mult_9_n156, mult_9_n104, mult_9_n103);
	xor gate_sum_13 (sum_13, mult_9_n105, mult_9_n157);
	xor gate_mult_9_n102 (mult_9_n102, mult_9_n596, mult_9_n567);
	and gate_mult_9_n101 (mult_9_n101, mult_9_n567, mult_9_n596);
	and gate_mult_9_n100 (mult_9_n100, mult_9_n156, mult_9_n102);
	or gate_mult_9_n155 (mult_9_n155, mult_9_n101, mult_9_n100);
	xor gate_sum_14 (sum_14, mult_9_n102, mult_9_n156);
	xor gate_mult_9_n99 (mult_9_n99, mult_9_n566, mult_9_n535);
	and gate_mult_9_n98 (mult_9_n98, mult_9_n535, mult_9_n566);
	and gate_mult_9_n97 (mult_9_n97, mult_9_n155, mult_9_n99);
	or gate_mult_9_n154 (mult_9_n154, mult_9_n98, mult_9_n97);
	xor gate_sum_15 (sum_15, mult_9_n99, mult_9_n155);
	xor gate_mult_9_n96 (mult_9_n96, mult_9_n534, mult_9_n500);
	and gate_mult_9_n95 (mult_9_n95, mult_9_n500, mult_9_n534);
	and gate_mult_9_n94 (mult_9_n94, mult_9_n154, mult_9_n96);
	or gate_mult_9_n153 (mult_9_n153, mult_9_n95, mult_9_n94);
	xor gate_sum_16 (sum_16, mult_9_n96, mult_9_n154);
	xor gate_mult_9_n93 (mult_9_n93, mult_9_n499, mult_9_n464);
	and gate_mult_9_n92 (mult_9_n92, mult_9_n464, mult_9_n499);
	and gate_mult_9_n91 (mult_9_n91, mult_9_n153, mult_9_n93);
	or gate_mult_9_n152 (mult_9_n152, mult_9_n92, mult_9_n91);
	xor gate_sum_17 (sum_17, mult_9_n93, mult_9_n153);
	xor gate_mult_9_n90 (mult_9_n90, mult_9_n463, mult_9_n427);
	and gate_mult_9_n89 (mult_9_n89, mult_9_n427, mult_9_n463);
	and gate_mult_9_n88 (mult_9_n88, mult_9_n152, mult_9_n90);
	or gate_mult_9_n151 (mult_9_n151, mult_9_n89, mult_9_n88);
	xor gate_sum_18 (sum_18, mult_9_n90, mult_9_n152);
	xor gate_mult_9_n87 (mult_9_n87, mult_9_n426, mult_9_n392);
	and gate_mult_9_n86 (mult_9_n86, mult_9_n392, mult_9_n426);
	and gate_mult_9_n85 (mult_9_n85, mult_9_n151, mult_9_n87);
	or gate_mult_9_n150 (mult_9_n150, mult_9_n86, mult_9_n85);
	xor gate_sum_19 (sum_19, mult_9_n87, mult_9_n151);
	xor gate_mult_9_n84 (mult_9_n84, mult_9_n391, mult_9_n360);
	and gate_mult_9_n83 (mult_9_n83, mult_9_n360, mult_9_n391);
	and gate_mult_9_n82 (mult_9_n82, mult_9_n150, mult_9_n84);
	or gate_mult_9_n149 (mult_9_n149, mult_9_n83, mult_9_n82);
	xor gate_sum_20 (sum_20, mult_9_n84, mult_9_n150);
	xor gate_mult_9_n81 (mult_9_n81, mult_9_n359, mult_9_n330);
	and gate_mult_9_n80 (mult_9_n80, mult_9_n330, mult_9_n359);
	and gate_mult_9_n79 (mult_9_n79, mult_9_n149, mult_9_n81);
	or gate_mult_9_n148 (mult_9_n148, mult_9_n80, mult_9_n79);
	xor gate_sum_21 (sum_21, mult_9_n81, mult_9_n149);
	xor gate_mult_9_n78 (mult_9_n78, mult_9_n329, mult_9_n303);
	and gate_mult_9_n77 (mult_9_n77, mult_9_n303, mult_9_n329);
	and gate_mult_9_n76 (mult_9_n76, mult_9_n148, mult_9_n78);
	or gate_mult_9_n147 (mult_9_n147, mult_9_n77, mult_9_n76);
	xor gate_sum_22 (sum_22, mult_9_n78, mult_9_n148);
	xor gate_mult_9_n75 (mult_9_n75, mult_9_n302, mult_9_n278);
	and gate_mult_9_n74 (mult_9_n74, mult_9_n278, mult_9_n302);
	and gate_mult_9_n73 (mult_9_n73, mult_9_n147, mult_9_n75);
	or gate_mult_9_n146 (mult_9_n146, mult_9_n74, mult_9_n73);
	xor gate_sum_23 (sum_23, mult_9_n75, mult_9_n147);
	xor gate_mult_9_n72 (mult_9_n72, mult_9_n277, mult_9_n256);
	and gate_mult_9_n71 (mult_9_n71, mult_9_n256, mult_9_n277);
	and gate_mult_9_n70 (mult_9_n70, mult_9_n146, mult_9_n72);
	or gate_mult_9_n145 (mult_9_n145, mult_9_n71, mult_9_n70);
	xor gate_sum_24 (sum_24, mult_9_n72, mult_9_n146);
	xor gate_mult_9_n69 (mult_9_n69, mult_9_n255, mult_9_n236);
	and gate_mult_9_n68 (mult_9_n68, mult_9_n236, mult_9_n255);
	and gate_mult_9_n67 (mult_9_n67, mult_9_n145, mult_9_n69);
	or gate_mult_9_n144 (mult_9_n144, mult_9_n68, mult_9_n67);
	xor gate_sum_25 (sum_25, mult_9_n69, mult_9_n145);
	xor gate_mult_9_n66 (mult_9_n66, mult_9_n219, mult_9_n235);
	and gate_mult_9_n65 (mult_9_n65, mult_9_n235, mult_9_n219);
	and gate_mult_9_n64 (mult_9_n64, mult_9_n144, mult_9_n66);
	or gate_mult_9_n143 (mult_9_n143, mult_9_n65, mult_9_n64);
	xor gate_sum_26 (sum_26, mult_9_n66, mult_9_n144);
	xor gate_mult_9_n63 (mult_9_n63, mult_9_n204, mult_9_n218);
	and gate_mult_9_n62 (mult_9_n62, mult_9_n218, mult_9_n204);
	and gate_mult_9_n61 (mult_9_n61, mult_9_n143, mult_9_n63);
	or gate_mult_9_n142 (mult_9_n142, mult_9_n62, mult_9_n61);
	xor gate_sum_27 (sum_27, mult_9_n63, mult_9_n143);
	xor gate_mult_9_n60 (mult_9_n60, mult_9_n203, mult_9_n192);
	and gate_mult_9_n59 (mult_9_n59, mult_9_n192, mult_9_n203);
	and gate_mult_9_n58 (mult_9_n58, mult_9_n142, mult_9_n60);
	or gate_mult_9_n141 (mult_9_n141, mult_9_n59, mult_9_n58);
	xor gate_sum_28 (sum_28, mult_9_n60, mult_9_n142);
	xor gate_mult_9_n57 (mult_9_n57, mult_9_n182, mult_9_n191);
	and gate_mult_9_n56 (mult_9_n56, mult_9_n191, mult_9_n182);
	and gate_mult_9_n55 (mult_9_n55, mult_9_n141, mult_9_n57);
	or gate_mult_9_n140 (mult_9_n140, mult_9_n56, mult_9_n55);
	xor gate_sum_29 (sum_29, mult_9_n57, mult_9_n141);
	xor gate_mult_9_n54 (mult_9_n54, mult_9_n175, mult_9_n181);
	and gate_mult_9_n53 (mult_9_n53, mult_9_n181, mult_9_n175);
	and gate_mult_9_n52 (mult_9_n52, mult_9_n140, mult_9_n54);
	or gate_mult_9_n139 (mult_9_n139, mult_9_n53, mult_9_n52);
	xor gate_sum_30 (sum_30, mult_9_n54, mult_9_n140);
	xor gate_mult_9_n51 (mult_9_n51, mult_9_n170, mult_9_n174);
	xor gate_sum_31 (sum_31, mult_9_n51, mult_9_n139);
	buf gate_mult_9_n49 (mult_9_n49, b_0);
	buf gate_mult_9_n48 (mult_9_n48, mult_9_n1387);
	buf gate_mult_9_n47 (mult_9_n47, mult_9_n1387);
	buf gate_mult_9_n46 (mult_9_n46, mult_9_n1396);
	buf gate_mult_9_n45 (mult_9_n45, mult_9_n1396);
	buf gate_mult_9_n43 (mult_9_n43, a_15);
	buf gate_mult_9_n42 (mult_9_n42, mult_9_n1388);
	buf gate_mult_9_n41 (mult_9_n41, mult_9_n1388);
	buf gate_mult_9_n40 (mult_9_n40, mult_9_n1397);
	buf gate_mult_9_n39 (mult_9_n39, mult_9_n1397);
	buf gate_mult_9_n37 (mult_9_n37, a_13);
	buf gate_mult_9_n36 (mult_9_n36, mult_9_n1389);
	buf gate_mult_9_n35 (mult_9_n35, mult_9_n1389);
	buf gate_mult_9_n34 (mult_9_n34, mult_9_n1398);
	buf gate_mult_9_n33 (mult_9_n33, mult_9_n1398);
	buf gate_mult_9_n31 (mult_9_n31, a_11);
	buf gate_mult_9_n30 (mult_9_n30, mult_9_n1390);
	buf gate_mult_9_n29 (mult_9_n29, mult_9_n1390);
	buf gate_mult_9_n28 (mult_9_n28, mult_9_n1399);
	buf gate_mult_9_n27 (mult_9_n27, mult_9_n1399);
	buf gate_mult_9_n25 (mult_9_n25, a_9);
	buf gate_mult_9_n24 (mult_9_n24, mult_9_n1391);
	buf gate_mult_9_n23 (mult_9_n23, mult_9_n1391);
	buf gate_mult_9_n22 (mult_9_n22, mult_9_n1400);
	buf gate_mult_9_n21 (mult_9_n21, mult_9_n1400);
	buf gate_mult_9_n19 (mult_9_n19, a_7);
	buf gate_mult_9_n18 (mult_9_n18, mult_9_n1392);
	buf gate_mult_9_n17 (mult_9_n17, mult_9_n1392);
	buf gate_mult_9_n16 (mult_9_n16, mult_9_n1401);
	buf gate_mult_9_n15 (mult_9_n15, mult_9_n1401);
	buf gate_mult_9_n13 (mult_9_n13, a_5);
	buf gate_mult_9_n12 (mult_9_n12, mult_9_n1393);
	buf gate_mult_9_n11 (mult_9_n11, mult_9_n1393);
	buf gate_mult_9_n10 (mult_9_n10, mult_9_n1402);
	buf gate_mult_9_n9 (mult_9_n9, mult_9_n1402);
	buf gate_mult_9_n7 (mult_9_n7, a_3);
	buf gate_mult_9_n6 (mult_9_n6, mult_9_n1394);
	buf gate_mult_9_n5 (mult_9_n5, mult_9_n1394);
	buf gate_mult_9_n4 (mult_9_n4, mult_9_n1403);
	buf gate_mult_9_n3 (mult_9_n3, mult_9_n1403);
	buf gate_mult_9_n1 (mult_9_n1, a_1);
endmodule

