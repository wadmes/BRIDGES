
module test ( a_0, a_1, a_2, a_3, a_4, a_5, a_6, a_7, b_0, b_1, b_2, b_3, b_4, b_5, b_6, b_7, 
  anoymous2_0, anoymous2_1, anoymous2_2, anoymous2_3, anoymous2_4, anoymous2_5, anoymous2_6, anoymous2_7, anoymous2_8, anoymous2_9, anoymous2_10, anoymous2_11, 
   anoymous2_12, anoymous2_13, anoymous2_14, anoymous2_15);
  
  input a_0;
  input a_1;
  input a_2;
  input a_3;
  input a_4;
  input a_5;
  input a_6;
  input a_7;

  input b_0;
  input b_1;
  input b_2;
  input b_3;
  input b_4;
  input b_5;
  input b_6;
  input b_7;
  
  output anoymous2_0;
  output anoymous2_1;
  output anoymous2_2;
  output anoymous2_3;
  output anoymous2_4;
  output anoymous2_5;
  output anoymous2_6;
  output anoymous2_7;
  output anoymous2_8;
  output anoymous2_9;
  output anoymous2_10;
  output anoymous2_11;
  output anoymous2_12;
  output anoymous2_13;
  output anoymous2_14;
  output anoymous2_15;
 

	not gate_anoymous_9_n321 (anoymous_9_n321, a_0);
	not gate_anoymous_9_n320 (anoymous_9_n320, a_1);
	not gate_anoymous_9_n319 (anoymous_9_n319, a_2);
	not gate_anoymous_9_n318 (anoymous_9_n318, a_3);
	not gate_anoymous_9_n317 (anoymous_9_n317, a_4);
	not gate_anoymous_9_n316 (anoymous_9_n316, a_5);
	not gate_anoymous_9_n315 (anoymous_9_n315, a_6);
	not gate_anoymous_9_n314 (anoymous_9_n314, a_7);
	not gate_anoymous_9_n313 (anoymous_9_n313, b_0);
	not gate_anoymous_9_n312 (anoymous_9_n312, b_1);
	not gate_anoymous_9_n311 (anoymous_9_n311, b_2);
	not gate_anoymous_9_n310 (anoymous_9_n310, b_3);
	not gate_anoymous_9_n309 (anoymous_9_n309, b_4);
	not gate_anoymous_9_n308 (anoymous_9_n308, b_5);
	not gate_anoymous_9_n307 (anoymous_9_n307, b_6);
	not gate_anoymous_9_n306 (anoymous_9_n306, b_7);
	nor gate_anoymous2_0 (anoymous2_0, anoymous_9_n321, anoymous_9_n313);
	nor gate_anoymous_9_n305 (anoymous_9_n305, anoymous_9_n321, anoymous_9_n312);
	nor gate_anoymous_9_n304 (anoymous_9_n304, anoymous_9_n321, anoymous_9_n311);
	nor gate_anoymous_9_n303 (anoymous_9_n303, anoymous_9_n321, anoymous_9_n310);
	nor gate_anoymous_9_n302 (anoymous_9_n302, anoymous_9_n321, anoymous_9_n309);
	nor gate_anoymous_9_n301 (anoymous_9_n301, anoymous_9_n321, anoymous_9_n308);
	nor gate_anoymous_9_n300 (anoymous_9_n300, anoymous_9_n321, anoymous_9_n307);
	nor gate_anoymous_9_n299 (anoymous_9_n299, anoymous_9_n321, anoymous_9_n306);
	nor gate_anoymous_9_n298 (anoymous_9_n298, anoymous_9_n320, anoymous_9_n313);
	nor gate_anoymous_9_n297 (anoymous_9_n297, anoymous_9_n320, anoymous_9_n312);
	nor gate_anoymous_9_n296 (anoymous_9_n296, anoymous_9_n320, anoymous_9_n311);
	nor gate_anoymous_9_n295 (anoymous_9_n295, anoymous_9_n320, anoymous_9_n310);
	nor gate_anoymous_9_n294 (anoymous_9_n294, anoymous_9_n320, anoymous_9_n309);
	nor gate_anoymous_9_n293 (anoymous_9_n293, anoymous_9_n320, anoymous_9_n308);
	nor gate_anoymous_9_n292 (anoymous_9_n292, anoymous_9_n320, anoymous_9_n307);
	nor gate_anoymous_9_n291 (anoymous_9_n291, anoymous_9_n320, anoymous_9_n306);
	nor gate_anoymous_9_n290 (anoymous_9_n290, anoymous_9_n319, anoymous_9_n313);
	nor gate_anoymous_9_n289 (anoymous_9_n289, anoymous_9_n319, anoymous_9_n312);
	nor gate_anoymous_9_n288 (anoymous_9_n288, anoymous_9_n319, anoymous_9_n311);
	nor gate_anoymous_9_n287 (anoymous_9_n287, anoymous_9_n319, anoymous_9_n310);
	nor gate_anoymous_9_n286 (anoymous_9_n286, anoymous_9_n319, anoymous_9_n309);
	nor gate_anoymous_9_n285 (anoymous_9_n285, anoymous_9_n319, anoymous_9_n308);
	nor gate_anoymous_9_n284 (anoymous_9_n284, anoymous_9_n319, anoymous_9_n307);
	nor gate_anoymous_9_n283 (anoymous_9_n283, anoymous_9_n319, anoymous_9_n306);
	nor gate_anoymous_9_n282 (anoymous_9_n282, anoymous_9_n318, anoymous_9_n313);
	nor gate_anoymous_9_n281 (anoymous_9_n281, anoymous_9_n318, anoymous_9_n312);
	nor gate_anoymous_9_n280 (anoymous_9_n280, anoymous_9_n318, anoymous_9_n311);
	nor gate_anoymous_9_n279 (anoymous_9_n279, anoymous_9_n318, anoymous_9_n310);
	nor gate_anoymous_9_n278 (anoymous_9_n278, anoymous_9_n318, anoymous_9_n309);
	nor gate_anoymous_9_n277 (anoymous_9_n277, anoymous_9_n318, anoymous_9_n308);
	nor gate_anoymous_9_n276 (anoymous_9_n276, anoymous_9_n318, anoymous_9_n307);
	nor gate_anoymous_9_n275 (anoymous_9_n275, anoymous_9_n318, anoymous_9_n306);
	nor gate_anoymous_9_n274 (anoymous_9_n274, anoymous_9_n317, anoymous_9_n313);
	nor gate_anoymous_9_n273 (anoymous_9_n273, anoymous_9_n317, anoymous_9_n312);
	nor gate_anoymous_9_n272 (anoymous_9_n272, anoymous_9_n317, anoymous_9_n311);
	nor gate_anoymous_9_n271 (anoymous_9_n271, anoymous_9_n317, anoymous_9_n310);
	nor gate_anoymous_9_n270 (anoymous_9_n270, anoymous_9_n317, anoymous_9_n309);
	nor gate_anoymous_9_n269 (anoymous_9_n269, anoymous_9_n317, anoymous_9_n308);
	nor gate_anoymous_9_n268 (anoymous_9_n268, anoymous_9_n317, anoymous_9_n307);
	nor gate_anoymous_9_n267 (anoymous_9_n267, anoymous_9_n317, anoymous_9_n306);
	nor gate_anoymous_9_n266 (anoymous_9_n266, anoymous_9_n316, anoymous_9_n313);
	nor gate_anoymous_9_n265 (anoymous_9_n265, anoymous_9_n316, anoymous_9_n312);
	nor gate_anoymous_9_n264 (anoymous_9_n264, anoymous_9_n316, anoymous_9_n311);
	nor gate_anoymous_9_n263 (anoymous_9_n263, anoymous_9_n316, anoymous_9_n310);
	nor gate_anoymous_9_n262 (anoymous_9_n262, anoymous_9_n316, anoymous_9_n309);
	nor gate_anoymous_9_n261 (anoymous_9_n261, anoymous_9_n316, anoymous_9_n308);
	nor gate_anoymous_9_n260 (anoymous_9_n260, anoymous_9_n316, anoymous_9_n307);
	nor gate_anoymous_9_n259 (anoymous_9_n259, anoymous_9_n316, anoymous_9_n306);
	nor gate_anoymous_9_n258 (anoymous_9_n258, anoymous_9_n315, anoymous_9_n313);
	nor gate_anoymous_9_n257 (anoymous_9_n257, anoymous_9_n315, anoymous_9_n312);
	nor gate_anoymous_9_n256 (anoymous_9_n256, anoymous_9_n315, anoymous_9_n311);
	nor gate_anoymous_9_n255 (anoymous_9_n255, anoymous_9_n315, anoymous_9_n310);
	nor gate_anoymous_9_n254 (anoymous_9_n254, anoymous_9_n315, anoymous_9_n309);
	nor gate_anoymous_9_n253 (anoymous_9_n253, anoymous_9_n315, anoymous_9_n308);
	nor gate_anoymous_9_n252 (anoymous_9_n252, anoymous_9_n315, anoymous_9_n307);
	nor gate_anoymous_9_n251 (anoymous_9_n251, anoymous_9_n315, anoymous_9_n306);
	nor gate_anoymous_9_n250 (anoymous_9_n250, anoymous_9_n314, anoymous_9_n313);
	nor gate_anoymous_9_n249 (anoymous_9_n249, anoymous_9_n314, anoymous_9_n312);
	nor gate_anoymous_9_n248 (anoymous_9_n248, anoymous_9_n314, anoymous_9_n311);
	nor gate_anoymous_9_n247 (anoymous_9_n247, anoymous_9_n314, anoymous_9_n310);
	nor gate_anoymous_9_n246 (anoymous_9_n246, anoymous_9_n314, anoymous_9_n309);
	nor gate_anoymous_9_n245 (anoymous_9_n245, anoymous_9_n314, anoymous_9_n308);
	nor gate_anoymous_9_n244 (anoymous_9_n244, anoymous_9_n314, anoymous_9_n307);
	nor gate_anoymous_9_n243 (anoymous_9_n243, anoymous_9_n314, anoymous_9_n306);
	and gate_anoymous_9_n241 (anoymous_9_n241, anoymous_9_n297, anoymous_9_n304);
	xor gate_anoymous_9_n242 (anoymous_9_n242, anoymous_9_n304, anoymous_9_n297);
	and gate_anoymous_9_n239 (anoymous_9_n239, anoymous_9_n282, anoymous_9_n289);
	xor gate_anoymous_9_n240 (anoymous_9_n240, anoymous_9_n289, anoymous_9_n282);
	xor gate_anoymous_9_n236 (anoymous_9_n236, anoymous_9_n303, anoymous_9_n296);
	and gate_anoymous_9_n235 (anoymous_9_n235, anoymous_9_n296, anoymous_9_n303);
	and gate_anoymous_9_n234 (anoymous_9_n234, anoymous_9_n236, anoymous_9_n241);
	or gate_anoymous_9_n237 (anoymous_9_n237, anoymous_9_n235, anoymous_9_n234);
	xor gate_anoymous_9_n238 (anoymous_9_n238, anoymous_9_n241, anoymous_9_n236);
	and gate_anoymous_9_n232 (anoymous_9_n232, anoymous_9_n274, anoymous_9_n281);
	xor gate_anoymous_9_n233 (anoymous_9_n233, anoymous_9_n281, anoymous_9_n274);
	xor gate_anoymous_9_n229 (anoymous_9_n229, anoymous_9_n302, anoymous_9_n295);
	and gate_anoymous_9_n228 (anoymous_9_n228, anoymous_9_n295, anoymous_9_n302);
	and gate_anoymous_9_n227 (anoymous_9_n227, anoymous_9_n229, anoymous_9_n288);
	or gate_anoymous_9_n230 (anoymous_9_n230, anoymous_9_n228, anoymous_9_n227);
	xor gate_anoymous_9_n231 (anoymous_9_n231, anoymous_9_n288, anoymous_9_n229);
	xor gate_anoymous_9_n224 (anoymous_9_n224, anoymous_9_n239, anoymous_9_n233);
	and gate_anoymous_9_n223 (anoymous_9_n223, anoymous_9_n233, anoymous_9_n239);
	and gate_anoymous_9_n222 (anoymous_9_n222, anoymous_9_n224, anoymous_9_n237);
	or gate_anoymous_9_n225 (anoymous_9_n225, anoymous_9_n223, anoymous_9_n222);
	xor gate_anoymous_9_n226 (anoymous_9_n226, anoymous_9_n237, anoymous_9_n224);
	and gate_anoymous_9_n220 (anoymous_9_n220, anoymous_9_n266, anoymous_9_n273);
	xor gate_anoymous_9_n221 (anoymous_9_n221, anoymous_9_n273, anoymous_9_n266);
	xor gate_anoymous_9_n217 (anoymous_9_n217, anoymous_9_n301, anoymous_9_n294);
	and gate_anoymous_9_n216 (anoymous_9_n216, anoymous_9_n294, anoymous_9_n301);
	and gate_anoymous_9_n215 (anoymous_9_n215, anoymous_9_n217, anoymous_9_n287);
	or gate_anoymous_9_n218 (anoymous_9_n218, anoymous_9_n216, anoymous_9_n215);
	xor gate_anoymous_9_n219 (anoymous_9_n219, anoymous_9_n287, anoymous_9_n217);
	xor gate_anoymous_9_n212 (anoymous_9_n212, anoymous_9_n280, anoymous_9_n232);
	and gate_anoymous_9_n211 (anoymous_9_n211, anoymous_9_n232, anoymous_9_n280);
	and gate_anoymous_9_n210 (anoymous_9_n210, anoymous_9_n212, anoymous_9_n221);
	or gate_anoymous_9_n213 (anoymous_9_n213, anoymous_9_n211, anoymous_9_n210);
	xor gate_anoymous_9_n214 (anoymous_9_n214, anoymous_9_n221, anoymous_9_n212);
	xor gate_anoymous_9_n207 (anoymous_9_n207, anoymous_9_n230, anoymous_9_n219);
	and gate_anoymous_9_n206 (anoymous_9_n206, anoymous_9_n219, anoymous_9_n230);
	and gate_anoymous_9_n205 (anoymous_9_n205, anoymous_9_n207, anoymous_9_n214);
	or gate_anoymous_9_n208 (anoymous_9_n208, anoymous_9_n206, anoymous_9_n205);
	xor gate_anoymous_9_n209 (anoymous_9_n209, anoymous_9_n214, anoymous_9_n207);
	and gate_anoymous_9_n203 (anoymous_9_n203, anoymous_9_n258, anoymous_9_n265);
	xor gate_anoymous_9_n204 (anoymous_9_n204, anoymous_9_n265, anoymous_9_n258);
	xor gate_anoymous_9_n200 (anoymous_9_n200, anoymous_9_n300, anoymous_9_n293);
	and gate_anoymous_9_n199 (anoymous_9_n199, anoymous_9_n293, anoymous_9_n300);
	and gate_anoymous_9_n198 (anoymous_9_n198, anoymous_9_n200, anoymous_9_n272);
	or gate_anoymous_9_n201 (anoymous_9_n201, anoymous_9_n199, anoymous_9_n198);
	xor gate_anoymous_9_n202 (anoymous_9_n202, anoymous_9_n272, anoymous_9_n200);
	xor gate_anoymous_9_n195 (anoymous_9_n195, anoymous_9_n286, anoymous_9_n279);
	and gate_anoymous_9_n194 (anoymous_9_n194, anoymous_9_n279, anoymous_9_n286);
	and gate_anoymous_9_n193 (anoymous_9_n193, anoymous_9_n195, anoymous_9_n220);
	or gate_anoymous_9_n196 (anoymous_9_n196, anoymous_9_n194, anoymous_9_n193);
	xor gate_anoymous_9_n197 (anoymous_9_n197, anoymous_9_n220, anoymous_9_n195);
	xor gate_anoymous_9_n190 (anoymous_9_n190, anoymous_9_n204, anoymous_9_n218);
	and gate_anoymous_9_n189 (anoymous_9_n189, anoymous_9_n218, anoymous_9_n204);
	and gate_anoymous_9_n188 (anoymous_9_n188, anoymous_9_n190, anoymous_9_n197);
	or gate_anoymous_9_n191 (anoymous_9_n191, anoymous_9_n189, anoymous_9_n188);
	xor gate_anoymous_9_n192 (anoymous_9_n192, anoymous_9_n197, anoymous_9_n190);
	xor gate_anoymous_9_n185 (anoymous_9_n185, anoymous_9_n202, anoymous_9_n213);
	and gate_anoymous_9_n184 (anoymous_9_n184, anoymous_9_n213, anoymous_9_n202);
	and gate_anoymous_9_n183 (anoymous_9_n183, anoymous_9_n208, anoymous_9_n185);
	or gate_anoymous_9_n186 (anoymous_9_n186, anoymous_9_n184, anoymous_9_n183);
	xor gate_anoymous_9_n187 (anoymous_9_n187, anoymous_9_n185, anoymous_9_n208);
	and gate_anoymous_9_n181 (anoymous_9_n181, anoymous_9_n250, anoymous_9_n257);
	xor gate_anoymous_9_n182 (anoymous_9_n182, anoymous_9_n257, anoymous_9_n250);
	xor gate_anoymous_9_n178 (anoymous_9_n178, anoymous_9_n299, anoymous_9_n292);
	and gate_anoymous_9_n177 (anoymous_9_n177, anoymous_9_n292, anoymous_9_n299);
	and gate_anoymous_9_n176 (anoymous_9_n176, anoymous_9_n178, anoymous_9_n271);
	or gate_anoymous_9_n179 (anoymous_9_n179, anoymous_9_n177, anoymous_9_n176);
	xor gate_anoymous_9_n180 (anoymous_9_n180, anoymous_9_n271, anoymous_9_n178);
	xor gate_anoymous_9_n173 (anoymous_9_n173, anoymous_9_n264, anoymous_9_n278);
	and gate_anoymous_9_n172 (anoymous_9_n172, anoymous_9_n278, anoymous_9_n264);
	and gate_anoymous_9_n171 (anoymous_9_n171, anoymous_9_n173, anoymous_9_n285);
	or gate_anoymous_9_n174 (anoymous_9_n174, anoymous_9_n172, anoymous_9_n171);
	xor gate_anoymous_9_n175 (anoymous_9_n175, anoymous_9_n285, anoymous_9_n173);
	xor gate_anoymous_9_n168 (anoymous_9_n168, anoymous_9_n203, anoymous_9_n182);
	and gate_anoymous_9_n167 (anoymous_9_n167, anoymous_9_n182, anoymous_9_n203);
	and gate_anoymous_9_n166 (anoymous_9_n166, anoymous_9_n168, anoymous_9_n201);
	or gate_anoymous_9_n169 (anoymous_9_n169, anoymous_9_n167, anoymous_9_n166);
	xor gate_anoymous_9_n170 (anoymous_9_n170, anoymous_9_n201, anoymous_9_n168);
	xor gate_anoymous_9_n163 (anoymous_9_n163, anoymous_9_n196, anoymous_9_n175);
	and gate_anoymous_9_n162 (anoymous_9_n162, anoymous_9_n175, anoymous_9_n196);
	and gate_anoymous_9_n161 (anoymous_9_n161, anoymous_9_n163, anoymous_9_n180);
	or gate_anoymous_9_n164 (anoymous_9_n164, anoymous_9_n162, anoymous_9_n161);
	xor gate_anoymous_9_n165 (anoymous_9_n165, anoymous_9_n180, anoymous_9_n163);
	xor gate_anoymous_9_n158 (anoymous_9_n158, anoymous_9_n170, anoymous_9_n191);
	and gate_anoymous_9_n157 (anoymous_9_n157, anoymous_9_n191, anoymous_9_n170);
	and gate_anoymous_9_n156 (anoymous_9_n156, anoymous_9_n158, anoymous_9_n165);
	or gate_anoymous_9_n159 (anoymous_9_n159, anoymous_9_n157, anoymous_9_n156);
	xor gate_anoymous_9_n160 (anoymous_9_n160, anoymous_9_n165, anoymous_9_n158);
	and gate_anoymous_9_n154 (anoymous_9_n154, anoymous_9_n249, anoymous_9_n256);
	xor gate_anoymous_9_n155 (anoymous_9_n155, anoymous_9_n256, anoymous_9_n249);
	xor gate_anoymous_9_n151 (anoymous_9_n151, anoymous_9_n270, anoymous_9_n277);
	and gate_anoymous_9_n150 (anoymous_9_n150, anoymous_9_n277, anoymous_9_n270);
	and gate_anoymous_9_n149 (anoymous_9_n149, anoymous_9_n151, anoymous_9_n263);
	or gate_anoymous_9_n152 (anoymous_9_n152, anoymous_9_n150, anoymous_9_n149);
	xor gate_anoymous_9_n153 (anoymous_9_n153, anoymous_9_n263, anoymous_9_n151);
	xor gate_anoymous_9_n146 (anoymous_9_n146, anoymous_9_n291, anoymous_9_n284);
	and gate_anoymous_9_n145 (anoymous_9_n145, anoymous_9_n284, anoymous_9_n291);
	and gate_anoymous_9_n144 (anoymous_9_n144, anoymous_9_n146, anoymous_9_n181);
	or gate_anoymous_9_n147 (anoymous_9_n147, anoymous_9_n145, anoymous_9_n144);
	xor gate_anoymous_9_n148 (anoymous_9_n148, anoymous_9_n181, anoymous_9_n146);
	xor gate_anoymous_9_n141 (anoymous_9_n141, anoymous_9_n155, anoymous_9_n179);
	and gate_anoymous_9_n140 (anoymous_9_n140, anoymous_9_n179, anoymous_9_n155);
	and gate_anoymous_9_n139 (anoymous_9_n139, anoymous_9_n141, anoymous_9_n174);
	or gate_anoymous_9_n142 (anoymous_9_n142, anoymous_9_n140, anoymous_9_n139);
	xor gate_anoymous_9_n143 (anoymous_9_n143, anoymous_9_n174, anoymous_9_n141);
	xor gate_anoymous_9_n136 (anoymous_9_n136, anoymous_9_n148, anoymous_9_n153);
	and gate_anoymous_9_n135 (anoymous_9_n135, anoymous_9_n153, anoymous_9_n148);
	and gate_anoymous_9_n134 (anoymous_9_n134, anoymous_9_n136, anoymous_9_n169);
	or gate_anoymous_9_n137 (anoymous_9_n137, anoymous_9_n135, anoymous_9_n134);
	xor gate_anoymous_9_n138 (anoymous_9_n138, anoymous_9_n169, anoymous_9_n136);
	xor gate_anoymous_9_n131 (anoymous_9_n131, anoymous_9_n164, anoymous_9_n143);
	and gate_anoymous_9_n130 (anoymous_9_n130, anoymous_9_n143, anoymous_9_n164);
	and gate_anoymous_9_n129 (anoymous_9_n129, anoymous_9_n131, anoymous_9_n138);
	or gate_anoymous_9_n132 (anoymous_9_n132, anoymous_9_n130, anoymous_9_n129);
	xor gate_anoymous_9_n133 (anoymous_9_n133, anoymous_9_n138, anoymous_9_n131);
	xor gate_anoymous_9_n126 (anoymous_9_n126, anoymous_9_n283, anoymous_9_n276);
	and gate_anoymous_9_n125 (anoymous_9_n125, anoymous_9_n276, anoymous_9_n283);
	and gate_anoymous_9_n124 (anoymous_9_n124, anoymous_9_n126, anoymous_9_n269);
	or gate_anoymous_9_n127 (anoymous_9_n127, anoymous_9_n125, anoymous_9_n124);
	xor gate_anoymous_9_n128 (anoymous_9_n128, anoymous_9_n269, anoymous_9_n126);
	xor gate_anoymous_9_n121 (anoymous_9_n121, anoymous_9_n262, anoymous_9_n255);
	and gate_anoymous_9_n120 (anoymous_9_n120, anoymous_9_n255, anoymous_9_n262);
	and gate_anoymous_9_n119 (anoymous_9_n119, anoymous_9_n121, anoymous_9_n248);
	or gate_anoymous_9_n122 (anoymous_9_n122, anoymous_9_n120, anoymous_9_n119);
	xor gate_anoymous_9_n123 (anoymous_9_n123, anoymous_9_n248, anoymous_9_n121);
	xor gate_anoymous_9_n116 (anoymous_9_n116, anoymous_9_n154, anoymous_9_n152);
	and gate_anoymous_9_n115 (anoymous_9_n115, anoymous_9_n152, anoymous_9_n154);
	and gate_anoymous_9_n114 (anoymous_9_n114, anoymous_9_n116, anoymous_9_n147);
	or gate_anoymous_9_n117 (anoymous_9_n117, anoymous_9_n115, anoymous_9_n114);
	xor gate_anoymous_9_n118 (anoymous_9_n118, anoymous_9_n147, anoymous_9_n116);
	xor gate_anoymous_9_n111 (anoymous_9_n111, anoymous_9_n123, anoymous_9_n128);
	and gate_anoymous_9_n110 (anoymous_9_n110, anoymous_9_n128, anoymous_9_n123);
	and gate_anoymous_9_n109 (anoymous_9_n109, anoymous_9_n142, anoymous_9_n111);
	or gate_anoymous_9_n112 (anoymous_9_n112, anoymous_9_n110, anoymous_9_n109);
	xor gate_anoymous_9_n113 (anoymous_9_n113, anoymous_9_n111, anoymous_9_n142);
	xor gate_anoymous_9_n106 (anoymous_9_n106, anoymous_9_n118, anoymous_9_n137);
	and gate_anoymous_9_n105 (anoymous_9_n105, anoymous_9_n137, anoymous_9_n118);
	and gate_anoymous_9_n104 (anoymous_9_n104, anoymous_9_n106, anoymous_9_n113);
	or gate_anoymous_9_n107 (anoymous_9_n107, anoymous_9_n105, anoymous_9_n104);
	xor gate_anoymous_9_n108 (anoymous_9_n108, anoymous_9_n113, anoymous_9_n106);
	xor gate_anoymous_9_n101 (anoymous_9_n101, anoymous_9_n275, anoymous_9_n268);
	and gate_anoymous_9_n100 (anoymous_9_n100, anoymous_9_n268, anoymous_9_n275);
	and gate_anoymous_9_n99 (anoymous_9_n99, anoymous_9_n101, anoymous_9_n261);
	or gate_anoymous_9_n102 (anoymous_9_n102, anoymous_9_n100, anoymous_9_n99);
	xor gate_anoymous_9_n103 (anoymous_9_n103, anoymous_9_n261, anoymous_9_n101);
	xor gate_anoymous_9_n96 (anoymous_9_n96, anoymous_9_n254, anoymous_9_n247);
	and gate_anoymous_9_n95 (anoymous_9_n95, anoymous_9_n247, anoymous_9_n254);
	and gate_anoymous_9_n94 (anoymous_9_n94, anoymous_9_n127, anoymous_9_n96);
	or gate_anoymous_9_n97 (anoymous_9_n97, anoymous_9_n95, anoymous_9_n94);
	xor gate_anoymous_9_n98 (anoymous_9_n98, anoymous_9_n96, anoymous_9_n127);
	xor gate_anoymous_9_n91 (anoymous_9_n91, anoymous_9_n122, anoymous_9_n103);
	and gate_anoymous_9_n90 (anoymous_9_n90, anoymous_9_n103, anoymous_9_n122);
	and gate_anoymous_9_n89 (anoymous_9_n89, anoymous_9_n91, anoymous_9_n98);
	or gate_anoymous_9_n92 (anoymous_9_n92, anoymous_9_n90, anoymous_9_n89);
	xor gate_anoymous_9_n93 (anoymous_9_n93, anoymous_9_n98, anoymous_9_n91);
	xor gate_anoymous_9_n86 (anoymous_9_n86, anoymous_9_n117, anoymous_9_n93);
	and gate_anoymous_9_n85 (anoymous_9_n85, anoymous_9_n93, anoymous_9_n117);
	and gate_anoymous_9_n84 (anoymous_9_n84, anoymous_9_n86, anoymous_9_n112);
	or gate_anoymous_9_n87 (anoymous_9_n87, anoymous_9_n85, anoymous_9_n84);
	xor gate_anoymous_9_n88 (anoymous_9_n88, anoymous_9_n112, anoymous_9_n86);
	xor gate_anoymous_9_n81 (anoymous_9_n81, anoymous_9_n267, anoymous_9_n260);
	and gate_anoymous_9_n80 (anoymous_9_n80, anoymous_9_n260, anoymous_9_n267);
	and gate_anoymous_9_n79 (anoymous_9_n79, anoymous_9_n81, anoymous_9_n253);
	or gate_anoymous_9_n82 (anoymous_9_n82, anoymous_9_n80, anoymous_9_n79);
	xor gate_anoymous_9_n83 (anoymous_9_n83, anoymous_9_n253, anoymous_9_n81);
	xor gate_anoymous_9_n76 (anoymous_9_n76, anoymous_9_n246, anoymous_9_n102);
	and gate_anoymous_9_n75 (anoymous_9_n75, anoymous_9_n102, anoymous_9_n246);
	and gate_anoymous_9_n74 (anoymous_9_n74, anoymous_9_n76, anoymous_9_n83);
	or gate_anoymous_9_n77 (anoymous_9_n77, anoymous_9_n75, anoymous_9_n74);
	xor gate_anoymous_9_n78 (anoymous_9_n78, anoymous_9_n83, anoymous_9_n76);
	xor gate_anoymous_9_n71 (anoymous_9_n71, anoymous_9_n97, anoymous_9_n92);
	and gate_anoymous_9_n70 (anoymous_9_n70, anoymous_9_n92, anoymous_9_n97);
	and gate_anoymous_9_n69 (anoymous_9_n69, anoymous_9_n71, anoymous_9_n78);
	or gate_anoymous_9_n72 (anoymous_9_n72, anoymous_9_n70, anoymous_9_n69);
	xor gate_anoymous_9_n73 (anoymous_9_n73, anoymous_9_n78, anoymous_9_n71);
	xor gate_anoymous_9_n66 (anoymous_9_n66, anoymous_9_n259, anoymous_9_n252);
	and gate_anoymous_9_n65 (anoymous_9_n65, anoymous_9_n252, anoymous_9_n259);
	and gate_anoymous_9_n64 (anoymous_9_n64, anoymous_9_n66, anoymous_9_n245);
	or gate_anoymous_9_n67 (anoymous_9_n67, anoymous_9_n65, anoymous_9_n64);
	xor gate_anoymous_9_n68 (anoymous_9_n68, anoymous_9_n245, anoymous_9_n66);
	xor gate_anoymous_9_n61 (anoymous_9_n61, anoymous_9_n82, anoymous_9_n68);
	and gate_anoymous_9_n60 (anoymous_9_n60, anoymous_9_n68, anoymous_9_n82);
	and gate_anoymous_9_n59 (anoymous_9_n59, anoymous_9_n77, anoymous_9_n61);
	or gate_anoymous_9_n62 (anoymous_9_n62, anoymous_9_n60, anoymous_9_n59);
	xor gate_anoymous_9_n63 (anoymous_9_n63, anoymous_9_n61, anoymous_9_n77);
	xor gate_anoymous_9_n56 (anoymous_9_n56, anoymous_9_n251, anoymous_9_n244);
	and gate_anoymous_9_n55 (anoymous_9_n55, anoymous_9_n244, anoymous_9_n251);
	and gate_anoymous_9_n54 (anoymous_9_n54, anoymous_9_n67, anoymous_9_n56);
	or gate_anoymous_9_n57 (anoymous_9_n57, anoymous_9_n55, anoymous_9_n54);
	xor gate_anoymous_9_n58 (anoymous_9_n58, anoymous_9_n56, anoymous_9_n67);
	and gate_anoymous_9_n53 (anoymous_9_n53, anoymous_9_n305, anoymous_9_n298);
	xor gate_anoymous2_1 (anoymous2_1, anoymous_9_n298, anoymous_9_n305);
	xor gate_anoymous_9_n39 (anoymous_9_n39, anoymous_9_n290, anoymous_9_n242);
	and gate_anoymous_9_n38 (anoymous_9_n38, anoymous_9_n242, anoymous_9_n290);
	and gate_anoymous_9_n37 (anoymous_9_n37, anoymous_9_n39, anoymous_9_n53);
	or gate_anoymous_9_n52 (anoymous_9_n52, anoymous_9_n38, anoymous_9_n37);
	xor gate_anoymous2_2 (anoymous2_2, anoymous_9_n53, anoymous_9_n39);
	xor gate_anoymous_9_n36 (anoymous_9_n36, anoymous_9_n240, anoymous_9_n238);
	and gate_anoymous_9_n35 (anoymous_9_n35, anoymous_9_n238, anoymous_9_n240);
	and gate_anoymous_9_n34 (anoymous_9_n34, anoymous_9_n36, anoymous_9_n52);
	or gate_anoymous_9_n51 (anoymous_9_n51, anoymous_9_n35, anoymous_9_n34);
	xor gate_anoymous2_3 (anoymous2_3, anoymous_9_n52, anoymous_9_n36);
	xor gate_anoymous_9_n33 (anoymous_9_n33, anoymous_9_n231, anoymous_9_n226);
	and gate_anoymous_9_n32 (anoymous_9_n32, anoymous_9_n226, anoymous_9_n231);
	and gate_anoymous_9_n31 (anoymous_9_n31, anoymous_9_n33, anoymous_9_n51);
	or gate_anoymous_9_n50 (anoymous_9_n50, anoymous_9_n32, anoymous_9_n31);
	xor gate_anoymous2_4 (anoymous2_4, anoymous_9_n51, anoymous_9_n33);
	xor gate_anoymous_9_n30 (anoymous_9_n30, anoymous_9_n225, anoymous_9_n209);
	and gate_anoymous_9_n29 (anoymous_9_n29, anoymous_9_n209, anoymous_9_n225);
	and gate_anoymous_9_n28 (anoymous_9_n28, anoymous_9_n30, anoymous_9_n50);
	or gate_anoymous_9_n49 (anoymous_9_n49, anoymous_9_n29, anoymous_9_n28);
	xor gate_anoymous2_5 (anoymous2_5, anoymous_9_n50, anoymous_9_n30);
	xor gate_anoymous_9_n27 (anoymous_9_n27, anoymous_9_n192, anoymous_9_n187);
	and gate_anoymous_9_n26 (anoymous_9_n26, anoymous_9_n187, anoymous_9_n192);
	and gate_anoymous_9_n25 (anoymous_9_n25, anoymous_9_n27, anoymous_9_n49);
	or gate_anoymous_9_n48 (anoymous_9_n48, anoymous_9_n26, anoymous_9_n25);
	xor gate_anoymous2_6 (anoymous2_6, anoymous_9_n49, anoymous_9_n27);
	xor gate_anoymous_9_n24 (anoymous_9_n24, anoymous_9_n186, anoymous_9_n160);
	and gate_anoymous_9_n23 (anoymous_9_n23, anoymous_9_n160, anoymous_9_n186);
	and gate_anoymous_9_n22 (anoymous_9_n22, anoymous_9_n48, anoymous_9_n24);
	or gate_anoymous_9_n47 (anoymous_9_n47, anoymous_9_n23, anoymous_9_n22);
	xor gate_anoymous2_7 (anoymous2_7, anoymous_9_n24, anoymous_9_n48);
	xor gate_anoymous_9_n21 (anoymous_9_n21, anoymous_9_n159, anoymous_9_n133);
	and gate_anoymous_9_n20 (anoymous_9_n20, anoymous_9_n133, anoymous_9_n159);
	and gate_anoymous_9_n19 (anoymous_9_n19, anoymous_9_n47, anoymous_9_n21);
	or gate_anoymous_9_n46 (anoymous_9_n46, anoymous_9_n20, anoymous_9_n19);
	xor gate_anoymous2_8 (anoymous2_8, anoymous_9_n21, anoymous_9_n47);
	xor gate_anoymous_9_n18 (anoymous_9_n18, anoymous_9_n132, anoymous_9_n108);
	and gate_anoymous_9_n17 (anoymous_9_n17, anoymous_9_n108, anoymous_9_n132);
	and gate_anoymous_9_n16 (anoymous_9_n16, anoymous_9_n46, anoymous_9_n18);
	or gate_anoymous_9_n45 (anoymous_9_n45, anoymous_9_n17, anoymous_9_n16);
	xor gate_anoymous2_9 (anoymous2_9, anoymous_9_n18, anoymous_9_n46);
	xor gate_anoymous_9_n15 (anoymous_9_n15, anoymous_9_n107, anoymous_9_n88);
	and gate_anoymous_9_n14 (anoymous_9_n14, anoymous_9_n88, anoymous_9_n107);
	and gate_anoymous_9_n13 (anoymous_9_n13, anoymous_9_n45, anoymous_9_n15);
	or gate_anoymous_9_n44 (anoymous_9_n44, anoymous_9_n14, anoymous_9_n13);
	xor gate_anoymous2_10 (anoymous2_10, anoymous_9_n15, anoymous_9_n45);
	xor gate_anoymous_9_n12 (anoymous_9_n12, anoymous_9_n87, anoymous_9_n73);
	and gate_anoymous_9_n11 (anoymous_9_n11, anoymous_9_n73, anoymous_9_n87);
	and gate_anoymous_9_n10 (anoymous_9_n10, anoymous_9_n44, anoymous_9_n12);
	or gate_anoymous_9_n43 (anoymous_9_n43, anoymous_9_n11, anoymous_9_n10);
	xor gate_anoymous2_11 (anoymous2_11, anoymous_9_n12, anoymous_9_n44);
	xor gate_anoymous_9_n9 (anoymous_9_n9, anoymous_9_n63, anoymous_9_n72);
	and gate_anoymous_9_n8 (anoymous_9_n8, anoymous_9_n72, anoymous_9_n63);
	and gate_anoymous_9_n7 (anoymous_9_n7, anoymous_9_n43, anoymous_9_n9);
	or gate_anoymous_9_n42 (anoymous_9_n42, anoymous_9_n8, anoymous_9_n7);
	xor gate_anoymous2_12 (anoymous2_12, anoymous_9_n9, anoymous_9_n43);
	xor gate_anoymous_9_n6 (anoymous_9_n6, anoymous_9_n58, anoymous_9_n62);
	and gate_anoymous_9_n5 (anoymous_9_n5, anoymous_9_n62, anoymous_9_n58);
	and gate_anoymous_9_n4 (anoymous_9_n4, anoymous_9_n42, anoymous_9_n6);
	or gate_anoymous_9_n41 (anoymous_9_n41, anoymous_9_n5, anoymous_9_n4);
	xor gate_anoymous2_13 (anoymous2_13, anoymous_9_n6, anoymous_9_n42);
	xor gate_anoymous_9_n3 (anoymous_9_n3, anoymous_9_n243, anoymous_9_n57);
	and gate_anoymous_9_n2 (anoymous_9_n2, anoymous_9_n57, anoymous_9_n243);
	and gate_anoymous_9_n1 (anoymous_9_n1, anoymous_9_n41, anoymous_9_n3);
	or gate_anoymous_9_n40 (anoymous_9_n40, anoymous_9_n2, anoymous_9_n1);
	xor gate_anoymous2_14 (anoymous2_14, anoymous_9_n3, anoymous_9_n41);
	buf gate_anoymous2_15 (anoymous2_15, anoymous_9_n40);
endmodule

